library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_sp_bits_1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_sp_bits_1 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"0B",X"AA",X"EA",X"00",X"BB",X"99",X"AE",X"00",X"BB",X"B9",X"A9",
		X"00",X"BA",X"B9",X"A9",X"99",X"AA",X"B9",X"9E",X"00",X"AA",X"BB",X"BB",X"00",X"AA",X"5B",X"BB",
		X"00",X"AA",X"55",X"B5",X"00",X"AA",X"66",X"55",X"0B",X"AA",X"5F",X"55",X"0B",X"55",X"FF",X"FF",
		X"0B",X"AA",X"5F",X"55",X"00",X"AA",X"55",X"55",X"00",X"AA",X"65",X"B5",X"00",X"AF",X"5B",X"BB",
		X"00",X"FF",X"BB",X"BB",X"99",X"AA",X"B9",X"99",X"00",X"B9",X"B9",X"A9",X"00",X"BB",X"B9",X"A9",
		X"00",X"BB",X"99",X"AE",X"00",X"0B",X"AA",X"EA",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"CA",X"00",X"00",X"00",
		X"AE",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"EB",X"AA",X"00",X"00",
		X"BB",X"BB",X"AA",X"00",X"BB",X"55",X"EB",X"AE",X"55",X"55",X"B5",X"55",X"5F",X"FF",X"FF",X"FF",
		X"55",X"55",X"B5",X"55",X"BB",X"55",X"EB",X"AE",X"BB",X"BB",X"AA",X"00",X"EB",X"AA",X"00",X"00",
		X"BE",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"AA",X"99",X"00",X"BB",X"BB",X"99",
		X"00",X"AA",X"BB",X"09",X"00",X"AA",X"BB",X"00",X"00",X"AA",X"9B",X"00",X"99",X"AA",X"BB",X"90",
		X"09",X"5A",X"BB",X"A9",X"00",X"A5",X"BB",X"A9",X"00",X"AA",X"BB",X"A9",X"00",X"A9",X"5B",X"A9",
		X"00",X"A9",X"55",X"99",X"00",X"F9",X"55",X"9B",X"00",X"A9",X"FA",X"BB",X"00",X"AA",X"FA",X"BB",
		X"00",X"A9",X"55",X"5B",X"00",X"B9",X"B5",X"55",X"00",X"BB",X"BB",X"55",X"00",X"AB",X"BB",X"FF",
		X"00",X"AA",X"A9",X"FF",X"00",X"0A",X"AA",X"55",X"00",X"00",X"AA",X"55",X"00",X"00",X"9A",X"BB",
		X"00",X"90",X"99",X"BB",X"00",X"09",X"99",X"BC",X"00",X"09",X"00",X"EB",X"00",X"00",X"00",X"BE",
		X"00",X"00",X"A0",X"AE",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"A0",X"00",X"00",
		X"B5",X"BA",X"00",X"00",X"BB",X"BB",X"00",X"00",X"AB",X"5B",X"00",X"00",X"AA",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"A0",X"00",X"00",X"AA",X"BA",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"AB",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"90",X"BB",X"00",X"00",X"90",X"BB",X"00",X"00",
		X"99",X"BB",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"AA",X"00",X"00",X"0B",X"AA",X"A0",X"00",
		X"0B",X"AA",X"BA",X"00",X"0B",X"5A",X"BA",X"00",X"0B",X"5A",X"B9",X"00",X"0B",X"55",X"BA",X"00",
		X"0B",X"BB",X"AA",X"90",X"0B",X"BB",X"AA",X"99",X"0B",X"B5",X"AA",X"99",X"0B",X"55",X"AA",X"09",
		X"0B",X"55",X"9A",X"09",X"00",X"55",X"9A",X"09",X"0A",X"B5",X"B9",X"99",X"00",X"B5",X"B9",X"99",
		X"00",X"BB",X"B9",X"00",X"00",X"BB",X"BB",X"00",X"00",X"9B",X"BB",X"00",X"99",X"9B",X"5B",X"00",
		X"99",X"99",X"5B",X"00",X"99",X"99",X"5B",X"00",X"99",X"99",X"F5",X"00",X"09",X"99",X"F5",X"00",
		X"09",X"99",X"F5",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"5F",X"00",X"00",X"99",X"BF",X"00",
		X"00",X"99",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"EB",X"A0",
		X"00",X"00",X"BE",X"A0",X"00",X"90",X"AB",X"A0",X"00",X"90",X"AA",X"AA",X"00",X"00",X"AA",X"CA",
		X"00",X"00",X"0A",X"AA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",
		X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"0E",X"5B",X"00",X"00",X"0B",X"5A",X"00",X"00",X"0B",X"5A",X"00",X"00",X"0B",X"5A",X"00",
		X"00",X"BB",X"5A",X"B0",X"00",X"BB",X"5A",X"B0",X"00",X"BB",X"5A",X"B0",X"00",X"AB",X"59",X"A0",
		X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"55",X"B0",X"00",X"AB",X"F5",X"A0",X"00",X"BB",X"FF",X"B0",
		X"00",X"AB",X"F5",X"A9",X"00",X"99",X"FF",X"99",X"00",X"99",X"AF",X"90",X"00",X"9A",X"AA",X"90",
		X"00",X"9A",X"AF",X"90",X"00",X"9A",X"FF",X"90",X"00",X"9A",X"F5",X"90",X"00",X"9A",X"FF",X"90",
		X"00",X"9A",X"F5",X"90",X"00",X"99",X"FF",X"99",X"00",X"AB",X"F5",X"A9",X"00",X"AE",X"55",X"A0",
		X"00",X"AB",X"F5",X"A0",X"00",X"AE",X"55",X"A0",X"00",X"AB",X"F5",X"A0",X"00",X"AE",X"55",X"A0",
		X"00",X"0A",X"55",X"00",X"00",X"0A",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"5A",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"05",X"F0",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"F5",X"50",X"00",X"00",X"F5",X"50",X"00",X"00",X"F5",X"F0",X"00",
		X"00",X"05",X"F3",X"00",X"00",X"00",X"F0",X"00",X"A0",X"05",X"05",X"3F",X"B0",X"05",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"F3",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"5F",X"F5",X"00",X"00",X"0F",X"50",X"00",X"00",X"F5",X"50",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"05",X"00",X"00",X"55",X"00",X"F0",X"00",X"50",X"05",X"00",X"00",X"00",X"00",X"05",
		X"00",X"50",X"00",X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"95",
		X"00",X"33",X"00",X"F5",X"00",X"30",X"00",X"55",X"00",X"59",X"00",X"95",X"00",X"55",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"74",X"00",X"00",X"00",
		X"74",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"71",X"00",X"00",X"60",X"66",X"00",X"00",X"F1",X"FF",
		X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"71",X"00",X"00",X"00",
		X"71",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"96",X"00",X"00",
		X"00",X"96",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"62",X"00",X"00",
		X"00",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"96",X"00",X"00",
		X"00",X"96",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"62",X"00",X"00",
		X"00",X"69",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"FA",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"FF",X"FA",X"00",X"00",X"FF",X"5A",X"00",X"00",X"F5",X"AE",X"00",
		X"00",X"F5",X"EE",X"00",X"00",X"F5",X"AE",X"00",X"00",X"F5",X"EE",X"00",X"00",X"F5",X"AE",X"00",
		X"00",X"0F",X"A5",X"00",X"00",X"0F",X"AF",X"00",X"00",X"0F",X"55",X"00",X"00",X"0F",X"55",X"00",
		X"00",X"0F",X"55",X"00",X"00",X"A0",X"5F",X"00",X"00",X"50",X"EF",X"00",X"00",X"50",X"E5",X"00",
		X"00",X"50",X"E5",X"00",X"00",X"05",X"5E",X"00",X"00",X"00",X"FE",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"0A",X"99",X"00",X"09",X"00",X"99",X"00",X"09",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"9D",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"9D",X"99",X"90",X"00",X"9D",X"99",X"90",
		X"00",X"9D",X"99",X"99",X"00",X"99",X"99",X"9D",X"00",X"99",X"99",X"9D",X"00",X"09",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9D",X"99",X"90",X"00",X"9D",X"99",X"90",
		X"00",X"9D",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"09",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"53",X"30",
		X"00",X"00",X"5E",X"30",X"00",X"00",X"55",X"30",X"00",X"00",X"E5",X"30",X"00",X"00",X"E5",X"00",
		X"00",X"00",X"53",X"00",X"00",X"03",X"55",X"00",X"00",X"05",X"F5",X"00",X"00",X"55",X"55",X"00",
		X"00",X"0F",X"F5",X"00",X"03",X"5E",X"05",X"00",X"FF",X"EE",X"F5",X"30",X"00",X"E5",X"F5",X"33",
		X"00",X"05",X"FF",X"E3",X"00",X"53",X"3F",X"E3",X"03",X"05",X"33",X"55",X"5F",X"55",X"E3",X"05",
		X"00",X"55",X"E5",X"50",X"00",X"55",X"35",X"33",X"00",X"FE",X"55",X"E3",X"00",X"0F",X"55",X"53",
		X"00",X"00",X"5E",X"50",X"00",X"00",X"5E",X"30",X"00",X"00",X"EE",X"30",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"50",X"00",X"05",X"53",X"E3",X"00",X"05",X"05",X"5E",X"00",X"55",X"55",X"5E",
		X"00",X"55",X"55",X"5E",X"00",X"55",X"55",X"E5",X"00",X"F5",X"55",X"E0",X"00",X"55",X"55",X"55",
		X"00",X"5F",X"55",X"55",X"00",X"F5",X"E5",X"E5",X"00",X"F5",X"5E",X"5E",X"00",X"05",X"55",X"5E",
		X"00",X"00",X"55",X"5E",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"05",X"55",X"F5",
		X"00",X"00",X"55",X"FF",X"00",X"EE",X"55",X"F5",X"00",X"E5",X"55",X"F5",X"00",X"55",X"55",X"3F",
		X"00",X"55",X"F5",X"30",X"00",X"55",X"E5",X"33",X"00",X"F5",X"53",X"5E",X"00",X"F5",X"E3",X"50",
		X"00",X"5F",X"E3",X"5E",X"00",X"55",X"EE",X"55",X"00",X"5F",X"5E",X"50",X"00",X"0F",X"5E",X"00",
		X"00",X"0F",X"5E",X"00",X"00",X"0F",X"E3",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"E9",X"99",X"00",X"00",X"BE",X"99",X"00",X"00",X"4B",X"99",X"00",X"00",X"74",X"EE",X"00",
		X"00",X"77",X"BE",X"90",X"00",X"34",X"5B",X"99",X"00",X"55",X"75",X"99",X"00",X"FF",X"99",X"EE",
		X"00",X"E5",X"95",X"BB",X"00",X"EE",X"99",X"99",X"00",X"F5",X"99",X"9F",X"55",X"55",X"95",X"F9",
		X"5F",X"5F",X"9F",X"F5",X"59",X"FF",X"9F",X"FF",X"59",X"FF",X"9F",X"FF",X"59",X"FF",X"FF",X"FF",
		X"0F",X"55",X"FF",X"FF",X"0F",X"55",X"FF",X"FF",X"EF",X"55",X"FF",X"F5",X"EF",X"75",X"FF",X"F5",
		X"EE",X"77",X"FF",X"F5",X"00",X"42",X"FF",X"F5",X"00",X"BB",X"55",X"F5",X"00",X"FF",X"99",X"F5",
		X"00",X"55",X"99",X"55",X"00",X"00",X"B9",X"55",X"00",X"00",X"FB",X"99",X"00",X"00",X"0F",X"99",
		X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"EA",X"90",X"00",X"00",X"EE",X"09",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"09",X"00",X"00",
		X"55",X"90",X"00",X"00",X"55",X"99",X"00",X"00",X"95",X"90",X"00",X"00",X"95",X"99",X"00",X"00",
		X"95",X"90",X"00",X"00",X"95",X"99",X"00",X"00",X"95",X"90",X"00",X"00",X"95",X"99",X"00",X"00",
		X"35",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"5E",X"00",X"00",X"00",X"54",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"3A",X"00",X"00",X"00",X"35",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"A9",X"00",
		X"00",X"49",X"A9",X"00",X"00",X"53",X"EA",X"00",X"00",X"55",X"EA",X"00",X"00",X"55",X"EA",X"00",
		X"00",X"59",X"EE",X"00",X"00",X"9F",X"4E",X"00",X"0A",X"FF",X"4E",X"00",X"0A",X"55",X"74",X"00",
		X"0A",X"F5",X"74",X"00",X"AA",X"55",X"54",X"00",X"0A",X"F5",X"57",X"00",X"00",X"55",X"57",X"00",
		X"00",X"F5",X"57",X"00",X"00",X"F5",X"55",X"00",X"00",X"5F",X"99",X"00",X"00",X"55",X"99",X"00",
		X"00",X"55",X"99",X"90",X"00",X"55",X"99",X"00",X"00",X"59",X"9F",X"90",X"00",X"99",X"FF",X"99",
		X"00",X"99",X"FF",X"90",X"00",X"99",X"FF",X"99",X"00",X"59",X"FF",X"A9",X"00",X"55",X"FF",X"A9",
		X"00",X"E5",X"FF",X"A9",X"00",X"E9",X"FF",X"AA",X"00",X"E9",X"FF",X"AA",X"00",X"E9",X"FF",X"EA",
		X"00",X"EE",X"FF",X"EA",X"00",X"EE",X"FF",X"EA",X"00",X"EE",X"FF",X"EE",X"00",X"AE",X"F9",X"9E",
		X"00",X"AE",X"99",X"9E",X"00",X"AE",X"F9",X"59",X"00",X"0A",X"55",X"54",X"00",X"0A",X"99",X"55",
		X"00",X"0A",X"95",X"53",X"00",X"00",X"99",X"53",X"00",X"00",X"99",X"54",X"00",X"00",X"99",X"54",
		X"00",X"00",X"53",X"44",X"00",X"00",X"55",X"EA",X"00",X"00",X"35",X"A3",X"00",X"00",X"33",X"35",
		X"00",X"00",X"33",X"35",X"00",X"00",X"43",X"35",X"00",X"00",X"AA",X"55",X"00",X"00",X"A1",X"99",
		X"00",X"00",X"A1",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"B0",X"F5",X"00",X"00",X"BB",X"F5",X"00",X"00",X"55",X"55",
		X"00",X"00",X"55",X"B5",X"00",X"00",X"55",X"5B",X"00",X"00",X"BB",X"55",X"00",X"00",X"BE",X"BB",
		X"00",X"00",X"BE",X"BB",X"00",X"00",X"5B",X"05",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",
		X"00",X"05",X"5B",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"5B",X"B0",X"00",X"5B",X"BB",X"B0",
		X"00",X"55",X"F5",X"B0",X"00",X"55",X"FF",X"B0",X"00",X"BB",X"5B",X"E0",X"00",X"55",X"B5",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"50",X"55",X"00",X"00",X"50",X"5B",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"BB",X"00",X"00",X"05",X"BB",X"00",
		X"00",X"55",X"BB",X"00",X"00",X"5F",X"BB",X"00",X"00",X"55",X"BB",X"00",X"00",X"5F",X"5F",X"00",
		X"00",X"5F",X"B5",X"00",X"00",X"55",X"5F",X"00",X"00",X"05",X"B5",X"00",X"00",X"05",X"5F",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"B0",X"BB",X"00",X"00",X"B0",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",
		X"09",X"99",X"99",X"05",X"AA",X"AA",X"99",X"FF",X"0A",X"EE",X"99",X"90",X"44",X"24",X"99",X"90",
		X"A7",X"37",X"99",X"99",X"AA",X"35",X"99",X"99",X"0A",X"33",X"99",X"AA",X"0A",X"53",X"9F",X"99",
		X"0A",X"55",X"5F",X"F9",X"09",X"55",X"5F",X"FF",X"09",X"55",X"FF",X"FF",X"09",X"59",X"FF",X"FF",
		X"09",X"59",X"F9",X"FF",X"0A",X"39",X"F9",X"FF",X"0A",X"39",X"F9",X"FF",X"0A",X"39",X"F9",X"F9",
		X"0A",X"39",X"99",X"99",X"AA",X"55",X"90",X"FF",X"A3",X"55",X"90",X"99",X"A7",X"77",X"33",X"F2",
		X"A4",X"2A",X"39",X"15",X"AE",X"EA",X"9F",X"EE",X"AA",X"9A",X"F3",X"AA",X"00",X"90",X"30",X"F3",
		X"00",X"00",X"39",X"09",X"00",X"00",X"9F",X"00",X"00",X"00",X"7F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"09",X"09",X"00",X"99",X"99",X"99",
		X"00",X"FF",X"99",X"05",X"00",X"EE",X"EE",X"EE",X"00",X"BB",X"BB",X"BB",X"0E",X"44",X"99",X"F5",
		X"0F",X"77",X"59",X"F9",X"5F",X"55",X"55",X"99",X"59",X"55",X"9F",X"55",X"59",X"FF",X"5F",X"FF",
		X"59",X"B5",X"FF",X"FF",X"5F",X"5E",X"FF",X"FF",X"5F",X"55",X"FF",X"FF",X"5F",X"55",X"FF",X"FF",
		X"5F",X"F5",X"FF",X"FF",X"5F",X"FF",X"FF",X"FF",X"5F",X"FF",X"FF",X"FF",X"59",X"FF",X"FF",X"FF",
		X"59",X"55",X"5F",X"FF",X"59",X"55",X"9F",X"55",X"5F",X"55",X"55",X"99",X"0F",X"77",X"F9",X"F9",
		X"0E",X"44",X"99",X"F5",X"00",X"BB",X"BB",X"BB",X"00",X"FF",X"FF",X"EF",X"00",X"FF",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"E9",X"90",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"90",X"00",X"00",
		X"44",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"B5",X"99",X"00",X"00",X"5B",X"99",X"00",X"00",
		X"35",X"59",X"00",X"00",X"93",X"59",X"00",X"00",X"93",X"59",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"93",X"59",X"00",X"00",X"93",X"59",X"00",X"00",X"35",X"59",X"00",X"00",
		X"55",X"90",X"00",X"00",X"55",X"09",X"00",X"00",X"FF",X"90",X"00",X"00",X"44",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"CC",X"CC",X"BC",X"00",X"EB",X"00",X"99",X"00",X"AA",X"BE",X"CC",X"99",X"AC",X"AA",X"BB",
		X"59",X"AA",X"EB",X"0B",X"59",X"BE",X"BE",X"C9",X"4C",X"EB",X"BB",X"BC",X"4C",X"BB",X"B5",X"EB",
		X"0C",X"BB",X"BB",X"BB",X"0C",X"EE",X"5B",X"BB",X"0C",X"5F",X"B5",X"BB",X"0C",X"BB",X"5B",X"BB",
		X"0C",X"BB",X"B5",X"BB",X"4C",X"BB",X"5B",X"BB",X"4C",X"BB",X"BF",X"69",X"50",X"66",X"FB",X"9B",
		X"50",X"BB",X"BB",X"BB",X"00",X"9C",X"6F",X"BB",X"00",X"EB",X"BB",X"CC",X"00",X"BE",X"00",X"99",
		X"00",X"CC",X"CC",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"97",X"99",X"99",X"00",X"77",X"9D",X"99",
		X"00",X"77",X"DD",X"99",X"00",X"00",X"DD",X"99",X"00",X"99",X"9A",X"E9",X"00",X"91",X"77",X"EE",
		X"9F",X"11",X"D7",X"EE",X"99",X"11",X"7D",X"EE",X"9F",X"1F",X"77",X"EE",X"99",X"1F",X"77",X"EE",
		X"00",X"01",X"77",X"EE",X"00",X"00",X"7D",X"E0",X"00",X"99",X"DD",X"00",X"00",X"77",X"7D",X"00",
		X"00",X"76",X"07",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"97",X"AA",X"AA",
		X"00",X"A3",X"9A",X"99",X"00",X"63",X"A9",X"99",X"00",X"66",X"9A",X"99",X"00",X"6F",X"A9",X"A3",
		X"00",X"66",X"99",X"3A",X"00",X"A9",X"A3",X"A0",X"00",X"99",X"A7",X"9F",X"00",X"FF",X"9A",X"9F",
		X"00",X"99",X"AA",X"9F",X"00",X"FF",X"AA",X"9F",X"00",X"99",X"99",X"9F",X"00",X"FF",X"55",X"9F",
		X"00",X"99",X"EA",X"9F",X"00",X"FF",X"AE",X"9F",X"00",X"99",X"EA",X"9F",X"00",X"FF",X"9E",X"9F",
		X"00",X"99",X"EA",X"9F",X"00",X"AA",X"EE",X"9F",X"00",X"66",X"99",X"E3",X"00",X"6F",X"A9",X"A3",
		X"00",X"66",X"EA",X"9E",X"00",X"6E",X"A9",X"99",X"00",X"EE",X"EA",X"99",X"00",X"9E",X"A9",X"99",
		X"00",X"35",X"D9",X"D9",X"00",X"D9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"A9",X"09",X"5E",X"90",
		X"99",X"99",X"EE",X"90",X"99",X"99",X"99",X"99",X"FF",X"FF",X"F9",X"99",X"99",X"99",X"99",X"44",
		X"9E",X"AA",X"57",X"AA",X"EA",X"AA",X"AA",X"55",X"EA",X"AA",X"AA",X"99",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"94",X"AA",X"AE",X"AA",X"49",X"AA",X"EE",X"EA",X"49",X"AA",X"E5",X"AA",X"A4",X"AA",X"E5",
		X"EA",X"A9",X"AA",X"E5",X"AE",X"94",X"AA",X"E5",X"EA",X"49",X"AA",X"EE",X"EE",X"49",X"AA",X"AE",
		X"EA",X"E4",X"AA",X"AA",X"5E",X"AE",X"AA",X"99",X"E5",X"EE",X"AE",X"55",X"9E",X"EE",X"55",X"AA",
		X"99",X"99",X"99",X"44",X"FF",X"FF",X"F9",X"99",X"99",X"99",X"99",X"99",X"99",X"D9",X"EE",X"90",
		X"D9",X"09",X"0E",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",
		X"00",X"EE",X"AA",X"AA",X"00",X"EE",X"99",X"EE",X"00",X"E5",X"93",X"55",X"00",X"99",X"3F",X"55",
		X"00",X"99",X"35",X"99",X"00",X"99",X"55",X"BA",X"09",X"94",X"FF",X"EE",X"09",X"43",X"FF",X"EE",
		X"09",X"49",X"FF",X"EE",X"09",X"94",X"FF",X"EE",X"09",X"AA",X"FF",X"EE",X"09",X"A4",X"FF",X"EE",
		X"09",X"49",X"FF",X"EE",X"09",X"49",X"F5",X"EE",X"09",X"47",X"55",X"EE",X"09",X"EE",X"55",X"B3",
		X"00",X"99",X"35",X"99",X"00",X"99",X"3F",X"55",X"00",X"EE",X"93",X"55",X"00",X"AA",X"99",X"EE",
		X"00",X"EE",X"EA",X"AE",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"A9",X"34",X"00",X"00",
		X"33",X"40",X"00",X"00",X"99",X"40",X"00",X"00",X"55",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"30",X"00",X"00",X"A5",X"90",X"00",X"00",
		X"55",X"A9",X"00",X"00",X"FF",X"A9",X"00",X"00",X"55",X"A9",X"00",X"00",X"55",X"A9",X"00",X"00",
		X"55",X"A9",X"00",X"00",X"A5",X"90",X"00",X"00",X"95",X"30",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"EE",X"40",X"00",X"00",
		X"99",X"40",X"00",X"00",X"A9",X"94",X"00",X"00",X"0E",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"90",X"90",X"99",X"00",X"09",X"09",X"99",X"00",X"99",X"90",X"22",
		X"00",X"99",X"99",X"22",X"92",X"33",X"99",X"22",X"FF",X"A3",X"99",X"22",X"F3",X"3A",X"22",X"22",
		X"F2",X"A3",X"92",X"22",X"09",X"99",X"29",X"22",X"93",X"33",X"29",X"22",X"92",X"95",X"29",X"22",
		X"99",X"55",X"29",X"22",X"9F",X"55",X"29",X"22",X"99",X"55",X"29",X"22",X"9F",X"55",X"29",X"22",
		X"99",X"99",X"29",X"22",X"9F",X"FF",X"29",X"22",X"99",X"FF",X"29",X"22",X"9F",X"FF",X"29",X"22",
		X"99",X"1F",X"29",X"22",X"92",X"1F",X"29",X"22",X"93",X"33",X"29",X"22",X"09",X"93",X"29",X"22",
		X"F2",X"A3",X"02",X"22",X"F2",X"3A",X"22",X"22",X"F2",X"A3",X"00",X"22",X"92",X"33",X"00",X"22",
		X"00",X"90",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"33",X"33",X"00",
		X"00",X"39",X"93",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"03",X"00",
		X"00",X"39",X"03",X"00",X"33",X"33",X"33",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"33",X"33",X"33",X"00",X"00",X"39",X"03",X"00",
		X"00",X"39",X"03",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"93",X"00",
		X"99",X"33",X"33",X"00",X"33",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"90",
		X"00",X"99",X"09",X"99",X"00",X"99",X"99",X"22",X"09",X"22",X"22",X"22",X"99",X"2D",X"22",X"22",
		X"9F",X"11",X"99",X"19",X"96",X"11",X"33",X"13",X"92",X"71",X"11",X"11",X"92",X"11",X"DD",X"7D",
		X"9F",X"11",X"D7",X"77",X"95",X"D1",X"77",X"77",X"95",X"4D",X"D7",X"77",X"95",X"44",X"75",X"77",
		X"95",X"44",X"77",X"77",X"95",X"44",X"75",X"77",X"95",X"57",X"F7",X"77",X"95",X"71",X"75",X"77",
		X"9F",X"11",X"F7",X"77",X"92",X"71",X"FF",X"FF",X"92",X"11",X"11",X"11",X"96",X"11",X"33",X"13",
		X"9F",X"77",X"99",X"19",X"99",X"F2",X"22",X"22",X"09",X"22",X"25",X"52",X"00",X"99",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"AA",X"00",X"00",X"00",X"11",X"90",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"90",X"00",X"00",X"92",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"92",X"00",X"00",X"00",X"11",X"90",X"00",X"00",
		X"11",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"09",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"90",X"90",X"90",X"90",X"00",
		X"00",X"05",X"00",X"50",X"00",X"05",X"53",X"E3",X"00",X"05",X"05",X"5E",X"50",X"55",X"55",X"5E",
		X"55",X"55",X"55",X"5E",X"55",X"55",X"55",X"E5",X"55",X"F5",X"55",X"E5",X"55",X"55",X"55",X"55",
		X"55",X"5F",X"55",X"55",X"55",X"F5",X"E5",X"E5",X"55",X"F5",X"5E",X"5E",X"55",X"55",X"55",X"5E",
		X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",
		X"55",X"55",X"55",X"FF",X"5F",X"EE",X"55",X"F5",X"5F",X"E5",X"55",X"F5",X"55",X"55",X"55",X"5F",
		X"5F",X"55",X"F5",X"55",X"55",X"55",X"E5",X"55",X"55",X"F5",X"55",X"5E",X"55",X"F5",X"E5",X"55",
		X"55",X"5F",X"E5",X"5E",X"55",X"55",X"EE",X"55",X"55",X"5F",X"5E",X"55",X"55",X"5F",X"5E",X"55",
		X"55",X"0F",X"55",X"55",X"05",X"0F",X"E3",X"53",X"05",X"00",X"00",X"53",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"30",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"93",X"33",X"00",
		X"00",X"00",X"39",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",
		X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",
		X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",
		X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",
		X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",
		X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",
		X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"19",X"90",X"00",
		X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"11",X"60",X"10",X"00",X"11",X"00",X"00",
		X"00",X"10",X"60",X"00",X"00",X"00",X"F1",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"91",X"00",
		X"00",X"01",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"19",X"00",X"00",X"19",X"19",X"90",
		X"00",X"19",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"91",X"00",X"00",X"11",X"91",X"00",X"00",X"11",X"91",X"09",
		X"00",X"11",X"91",X"91",X"00",X"99",X"9F",X"11",X"00",X"99",X"00",X"11",X"00",X"99",X"F0",X"10",
		X"00",X"99",X"6F",X"00",X"00",X"FF",X"66",X"00",X"00",X"90",X"66",X"11",X"01",X"11",X"6F",X"11",
		X"01",X"11",X"66",X"11",X"00",X"11",X"06",X"11",X"00",X"19",X"F9",X"11",X"00",X"90",X"0D",X"99",
		X"00",X"00",X"D1",X"00",X"00",X"00",X"11",X"10",X"00",X"09",X"11",X"10",X"00",X"91",X"11",X"11",
		X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"91",X"00",X"02",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"90",X"10",X"00",
		X"00",X"19",X"11",X"00",X"00",X"19",X"00",X"00",X"00",X"11",X"10",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"44",X"44",X"00",X"00",X"00",X"11",X"66",X"60",
		X"00",X"11",X"00",X"00",X"00",X"44",X"00",X"99",X"00",X"99",X"66",X"96",X"00",X"00",X"00",X"06",
		X"00",X"01",X"66",X"66",X"00",X"41",X"60",X"06",X"00",X"11",X"00",X"06",X"00",X"41",X"00",X"06",
		X"00",X"01",X"11",X"06",X"00",X"90",X"11",X"00",X"00",X"00",X"40",X"11",X"00",X"00",X"40",X"10",
		X"00",X"00",X"04",X"11",X"00",X"00",X"04",X"40",X"00",X"00",X"00",X"44",X"00",X"04",X"00",X"44",
		X"00",X"04",X"00",X"44",X"00",X"04",X"00",X"04",X"00",X"04",X"04",X"00",X"00",X"04",X"44",X"00",
		X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"10",X"09",X"00",X"00",X"41",X"99",X"09",X"00",X"41",X"44",X"09",X"00",X"91",X"11",X"09",X"00",
		X"91",X"09",X"01",X"09",X"55",X"10",X"11",X"90",X"51",X"00",X"41",X"04",X"55",X"00",X"11",X"44",
		X"59",X"00",X"44",X"14",X"50",X"00",X"66",X"40",X"50",X"00",X"60",X"00",X"55",X"66",X"01",X"00",
		X"50",X"60",X"01",X"00",X"5F",X"66",X"66",X"90",X"F6",X"00",X"66",X"49",X"F0",X"06",X"11",X"11",
		X"F0",X"00",X"00",X"44",X"5F",X"00",X"60",X"44",X"99",X"90",X"06",X"00",X"99",X"FF",X"00",X"00",
		X"06",X"F0",X"11",X"00",X"00",X"00",X"10",X"10",X"60",X"00",X"10",X"00",X"00",X"01",X"00",X"00",
		X"00",X"11",X"11",X"10",X"00",X"11",X"00",X"00",X"10",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"39",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"11",X"00",X"00",X"90",X"13",X"00",
		X"00",X"39",X"33",X"00",X"00",X"33",X"36",X"33",X"00",X"33",X"61",X"39",X"00",X"33",X"13",X"30",
		X"00",X"03",X"41",X"00",X"00",X"33",X"64",X"90",X"00",X"03",X"FF",X"00",X"00",X"36",X"F4",X"00",
		X"00",X"66",X"66",X"00",X"00",X"64",X"46",X"00",X"00",X"63",X"46",X"30",X"00",X"33",X"41",X"33",
		X"00",X"33",X"61",X"39",X"00",X"33",X"61",X"33",X"00",X"61",X"61",X"03",X"00",X"61",X"66",X"03",
		X"00",X"33",X"36",X"00",X"00",X"30",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"90",X"90",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"90",X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"90",
		X"00",X"39",X"66",X"99",X"60",X"36",X"66",X"99",X"66",X"93",X"66",X"99",X"00",X"36",X"61",X"96",
		X"00",X"93",X"11",X"69",X"00",X"13",X"16",X"31",X"01",X"66",X"FF",X"19",X"66",X"F1",X"FF",X"99",
		X"06",X"FF",X"FF",X"99",X"00",X"61",X"F1",X"99",X"00",X"66",X"46",X"99",X"00",X"44",X"F6",X"99",
		X"00",X"33",X"1F",X"90",X"00",X"66",X"1F",X"90",X"00",X"66",X"11",X"99",X"00",X"6F",X"69",X"99",
		X"09",X"66",X"69",X"99",X"99",X"66",X"69",X"69",X"99",X"66",X"69",X"99",X"90",X"69",X"69",X"66",
		X"00",X"66",X"99",X"99",X"00",X"00",X"96",X"99",X"00",X"00",X"96",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"09",X"09",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"93",X"99",X"90",
		X"00",X"93",X"99",X"39",X"00",X"99",X"39",X"39",X"00",X"99",X"39",X"93",X"00",X"99",X"91",X"39",
		X"00",X"96",X"61",X"93",X"00",X"93",X"61",X"39",X"00",X"93",X"33",X"93",X"00",X"96",X"19",X"99",
		X"00",X"30",X"11",X"99",X"00",X"00",X"31",X"19",X"00",X"63",X"99",X"99",X"00",X"16",X"61",X"99",
		X"00",X"33",X"19",X"99",X"00",X"63",X"19",X"39",X"00",X"33",X"11",X"39",X"00",X"44",X"61",X"99",
		X"00",X"36",X"99",X"39",X"00",X"33",X"96",X"30",X"00",X"09",X"16",X"99",X"00",X"33",X"99",X"99",
		X"00",X"33",X"99",X"33",X"09",X"31",X"91",X"13",X"09",X"33",X"99",X"61",X"09",X"99",X"99",X"69",
		X"00",X"33",X"99",X"99",X"00",X"09",X"61",X"99",X"00",X"00",X"33",X"99",X"00",X"00",X"39",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"39",X"99",X"00",
		X"00",X"39",X"13",X"30",X"00",X"33",X"33",X"00",X"00",X"93",X"99",X"00",X"00",X"19",X"99",X"00",
		X"00",X"16",X"99",X"00",X"00",X"66",X"63",X"90",X"00",X"33",X"33",X"93",X"00",X"31",X"33",X"33",
		X"00",X"91",X"39",X"93",X"00",X"13",X"33",X"39",X"00",X"39",X"19",X"39",X"00",X"30",X"99",X"00",
		X"00",X"31",X"99",X"33",X"00",X"11",X"33",X"99",X"03",X"41",X"33",X"39",X"00",X"06",X"99",X"39",
		X"00",X"09",X"13",X"33",X"00",X"19",X"93",X"39",X"09",X"11",X"99",X"90",X"00",X"99",X"39",X"39",
		X"00",X"90",X"93",X"33",X"00",X"99",X"11",X"33",X"00",X"90",X"66",X"39",X"00",X"30",X"16",X"39",
		X"00",X"99",X"99",X"39",X"00",X"00",X"39",X"99",X"00",X"90",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"39",X"00",
		X"00",X"03",X"99",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"93",X"39",X"00",X"33",X"93",X"30",X"00",X"33",X"39",X"93",
		X"00",X"33",X"39",X"93",X"00",X"39",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"93",X"93",X"00",
		X"00",X"93",X"39",X"00",X"00",X"33",X"39",X"00",X"00",X"39",X"39",X"90",X"00",X"99",X"39",X"39",
		X"00",X"90",X"99",X"39",X"00",X"00",X"93",X"30",X"00",X"00",X"30",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"50",X"F0",X"39",X"00",X"55",X"F0",X"90",
		X"00",X"55",X"3F",X"00",X"00",X"35",X"93",X"93",X"00",X"3F",X"99",X"30",X"00",X"33",X"99",X"30",
		X"00",X"5F",X"33",X"33",X"00",X"5F",X"93",X"33",X"00",X"93",X"33",X"53",X"00",X"35",X"93",X"93",
		X"00",X"55",X"33",X"90",X"00",X"55",X"93",X"33",X"00",X"55",X"33",X"33",X"00",X"99",X"99",X"33",
		X"00",X"55",X"99",X"53",X"00",X"55",X"33",X"30",X"00",X"53",X"FF",X"35",X"00",X"05",X"F0",X"33",
		X"00",X"00",X"F0",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"07",X"FF",X"04",
		X"00",X"07",X"FF",X"60",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"07",X"FF",X"06",
		X"00",X"77",X"FF",X"10",X"00",X"07",X"AA",X"60",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"7F",X"FF",X"04",
		X"00",X"77",X"FF",X"40",X"00",X"7F",X"AA",X"60",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"FF",X"06",
		X"00",X"FF",X"FF",X"61",X"00",X"FF",X"AA",X"10",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"FF",X"AA",X"00",X"07",X"FF",X"55",X"00",X"77",X"FF",X"FF",X"06",
		X"77",X"FF",X"FF",X"61",X"00",X"FF",X"AA",X"22",X"00",X"00",X"AA",X"22",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"FF",X"AA",X"00",X"07",X"FF",X"55",X"40",X"77",X"FF",X"FF",X"06",
		X"77",X"FF",X"FF",X"46",X"00",X"FF",X"AA",X"22",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"69",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"69",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"96",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"40",X"50",X"00",X"00",X"44",X"50",
		X"00",X"00",X"64",X"50",X"00",X"0F",X"44",X"00",X"00",X"00",X"64",X"00",X"00",X"0F",X"64",X"00",
		X"00",X"00",X"66",X"00",X"00",X"44",X"FF",X"30",X"00",X"33",X"FF",X"30",X"00",X"00",X"FF",X"50",
		X"00",X"00",X"66",X"00",X"00",X"03",X"66",X"40",X"00",X"0F",X"46",X"50",X"00",X"0F",X"44",X"00",
		X"00",X"0F",X"F4",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"5F",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"55",X"00",X"50",X"00",X"55",X"F0",X"50",
		X"00",X"55",X"45",X"50",X"00",X"5F",X"4F",X"00",X"00",X"55",X"64",X"00",X"00",X"5F",X"64",X"00",
		X"00",X"50",X"66",X"00",X"00",X"44",X"FF",X"35",X"00",X"33",X"FF",X"35",X"00",X"33",X"FF",X"55",
		X"00",X"E5",X"66",X"5F",X"00",X"53",X"6F",X"50",X"00",X"0F",X"4F",X"50",X"00",X"0F",X"F4",X"00",
		X"00",X"0F",X"FF",X"F0",X"00",X"00",X"54",X"00",X"00",X"00",X"5F",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"30",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"03",X"00",X"00",X"00",X"00",X"00",X"5E",X"00",X"00",X"55",X"0E",X"5E",X"00",X"55",X"55",X"5E",
		X"00",X"55",X"55",X"5E",X"00",X"5F",X"F3",X"50",X"00",X"5F",X"FF",X"50",X"00",X"5F",X"55",X"00",
		X"00",X"5F",X"55",X"33",X"00",X"55",X"5F",X"35",X"00",X"33",X"3F",X"35",X"00",X"33",X"FF",X"55",
		X"00",X"E5",X"FF",X"5F",X"00",X"53",X"55",X"55",X"00",X"FF",X"FF",X"55",X"00",X"5F",X"5F",X"55",
		X"00",X"FF",X"5F",X"F5",X"00",X"F5",X"55",X"E5",X"00",X"FF",X"5F",X"55",X"00",X"3F",X"55",X"50",
		X"00",X"5F",X"3F",X"50",X"00",X"5F",X"FF",X"05",X"00",X"EF",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"30",X"00",X"00",X"EE",X"00",X"00",X"00",X"E5",X"EE",X"00",X"00",X"E5",X"E5",X"00",
		X"00",X"55",X"5F",X"00",X"00",X"5F",X"FF",X"E0",X"00",X"5F",X"55",X"E0",X"00",X"55",X"EE",X"EE",
		X"00",X"55",X"F3",X"5E",X"00",X"5F",X"F5",X"5E",X"00",X"EE",X"FE",X"5E",X"00",X"35",X"FE",X"5E",
		X"00",X"EF",X"5F",X"5E",X"00",X"E3",X"5F",X"EE",X"00",X"FF",X"5F",X"E0",X"00",X"FE",X"F5",X"E0",
		X"00",X"F3",X"3F",X"00",X"00",X"35",X"3F",X"30",X"00",X"55",X"55",X"33",X"00",X"53",X"F3",X"50",
		X"00",X"53",X"35",X"E3",X"00",X"53",X"35",X"E3",X"00",X"55",X"FF",X"E0",X"00",X"F5",X"3F",X"E0",
		X"00",X"55",X"EE",X"00",X"00",X"FF",X"33",X"00",X"00",X"5F",X"0E",X"00",X"00",X"E5",X"03",X"33",
		X"00",X"E5",X"00",X"35",X"00",X"EE",X"00",X"33",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"64",X"64",X"00",
		X"00",X"46",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"44",X"00",
		X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"64",X"00",
		X"00",X"10",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"66",X"10",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"00",X"00",X"00",X"64",X"60",X"00",
		X"00",X"A6",X"16",X"00",X"00",X"66",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"16",X"06",X"40",
		X"00",X"66",X"66",X"46",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"64",X"60",X"00",X"00",X"11",X"06",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"60",X"40",
		X"00",X"16",X"06",X"00",X"00",X"10",X"00",X"00",X"00",X"66",X"01",X"00",X"00",X"A6",X"06",X"00",
		X"00",X"64",X"60",X"00",X"00",X"46",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"66",X"00",X"00",
		X"00",X"60",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"11",X"64",X"00",X"00",X"66",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"66",X"44",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"06",X"06",X"00",X"46",X"60",X"00",
		X"00",X"64",X"64",X"00",X"00",X"11",X"00",X"00",X"00",X"44",X"A0",X"00",X"00",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",X"00",X"90",X"00",X"91",X"09",X"09",
		X"00",X"11",X"90",X"90",X"00",X"11",X"99",X"09",X"00",X"11",X"99",X"90",X"00",X"91",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"7D",X"92",X"00",X"00",X"7D",X"22",X"00",X"06",X"7A",X"22",
		X"00",X"07",X"7A",X"29",X"00",X"77",X"AA",X"90",X"00",X"77",X"AD",X"09",X"00",X"00",X"DD",X"90",
		X"00",X"00",X"DA",X"49",X"00",X"00",X"DA",X"59",X"00",X"00",X"DD",X"59",X"00",X"00",X"DD",X"99",
		X"00",X"00",X"6D",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"55",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E9",X"00",X"00",X"DD",X"E9",
		X"00",X"00",X"77",X"E9",X"00",X"07",X"77",X"9A",X"00",X"07",X"7D",X"AD",X"00",X"70",X"D7",X"DD",
		X"00",X"17",X"7D",X"DD",X"00",X"10",X"7D",X"D9",X"00",X"90",X"2D",X"90",X"00",X"99",X"27",X"00",
		X"00",X"99",X"29",X"00",X"00",X"95",X"79",X"00",X"00",X"4E",X"79",X"00",X"00",X"6E",X"69",X"00",
		X"00",X"66",X"90",X"00",X"00",X"96",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"99",X"99",X"00",X"BF",X"96",X"99",X"00",X"00",X"64",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"99",X"99",X"04",X"0B",X"AF",X"4A",X"00",X"BB",X"FF",X"AE",X"00",X"BB",X"56",X"EE",
		X"00",X"00",X"56",X"E9",X"94",X"00",X"55",X"11",X"00",X"40",X"51",X"B0",X"00",X"F4",X"5F",X"11",
		X"00",X"F4",X"1F",X"11",X"00",X"FF",X"FF",X"FF",X"0B",X"AF",X"FF",X"55",X"00",X"FF",X"FF",X"1F",
		X"0A",X"F0",X"FF",X"55",X"66",X"00",X"FF",X"05",X"00",X"6F",X"65",X"05",X"00",X"66",X"51",X"BB",
		X"00",X"66",X"00",X"0B",X"99",X"66",X"FF",X"99",X"0F",X"06",X"BF",X"FF",X"00",X"06",X"6F",X"00",
		X"00",X"66",X"66",X"A0",X"00",X"BB",X"66",X"EA",X"00",X"B0",X"99",X"19",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"10",X"00",X"00",X"01",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"F1",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"11",X"00",X"00",X"40",X"0A",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"44",X"01",X"00",X"10",X"00",X"11",
		X"00",X"00",X"66",X"41",X"00",X"00",X"06",X"41",X"00",X"00",X"06",X"F1",X"00",X"00",X"11",X"F1",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"06",X"10",X"00",X"00",X"06",X"10",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"00",X"EB",X"00",X"69",X"00",X"03",X"00",X"40",X"66",X"0E",X"00",
		X"11",X"6E",X"00",X"00",X"11",X"0E",X"00",X"00",X"16",X"0E",X"00",X"00",X"11",X"00",X"11",X"00",
		X"16",X"66",X"10",X"00",X"66",X"00",X"10",X"00",X"16",X"11",X"00",X"00",X"16",X"00",X"00",X"00",
		X"66",X"16",X"00",X"BB",X"F6",X"66",X"00",X"E0",X"66",X"6B",X"BB",X"00",X"FF",X"56",X"11",X"EE",
		X"00",X"00",X"66",X"FF",X"00",X"00",X"01",X"01",X"00",X"00",X"11",X"01",X"00",X"00",X"00",X"FF",
		X"00",X"01",X"11",X"6F",X"00",X"01",X"01",X"66",X"00",X"00",X"01",X"66",X"00",X"00",X"10",X"66",
		X"00",X"00",X"66",X"61",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"B0",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"44",X"EE",X"00",X"F6",X"44",X"BB",X"00",X"66",X"66",X"66",X"0B",X"66",X"66",X"00",X"00",
		X"66",X"11",X"11",X"11",X"66",X"44",X"01",X"00",X"66",X"44",X"11",X"00",X"66",X"11",X"00",X"00",
		X"66",X"66",X"00",X"00",X"66",X"11",X"60",X"00",X"66",X"01",X"06",X"00",X"16",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"11",X"00",X"10",X"00",X"11",X"06",X"11",X"00",X"11",X"00",X"00",X"00",
		X"11",X"01",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"61",X"00",X"00",X"66",X"61",
		X"00",X"00",X"10",X"66",X"00",X"00",X"01",X"66",X"00",X"01",X"01",X"66",X"00",X"01",X"11",X"6F",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"11",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"66",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"01",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"06",X"11",X"00",X"11",X"00",X"10",X"00",X"16",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"66",X"01",X"06",X"00",X"66",X"11",X"60",X"00",X"66",X"66",X"00",X"00",
		X"66",X"11",X"00",X"00",X"66",X"44",X"11",X"00",X"66",X"44",X"01",X"00",X"61",X"11",X"11",X"11",
		X"11",X"66",X"00",X"00",X"16",X"66",X"66",X"0B",X"F6",X"44",X"BB",X"00",X"F6",X"44",X"EE",X"00",
		X"00",X"00",X"11",X"F1",X"00",X"00",X"06",X"F1",X"00",X"00",X"06",X"41",X"00",X"00",X"66",X"41",
		X"00",X"10",X"00",X"11",X"00",X"00",X"44",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"40",X"0A",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"1F",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"F1",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"56",X"11",X"EE",X"66",X"6B",X"00",X"00",X"F6",X"66",X"00",X"00",X"66",X"16",X"00",X"00",
		X"16",X"10",X"00",X"00",X"16",X"11",X"60",X"00",X"56",X"00",X"10",X"00",X"56",X"66",X"16",X"00",
		X"51",X"10",X"11",X"00",X"66",X"11",X"10",X"00",X"16",X"0E",X"10",X"00",X"11",X"6E",X"10",X"00",
		X"40",X"66",X"0E",X"00",X"69",X"00",X"03",X"00",X"66",X"00",X"EB",X"00",X"66",X"00",X"00",X"00",
		X"06",X"11",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"06",X"00",X"00",
		X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"04",X"01",X"00",X"00",X"00",X"11",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"41",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"43",X"66",X"00",X"00",
		X"11",X"60",X"00",X"00",X"16",X"33",X"00",X"00",X"30",X"11",X"10",X"00",X"33",X"33",X"00",X"00",
		X"00",X"66",X"16",X"00",X"30",X"33",X"10",X"00",X"33",X"03",X"60",X"00",X"03",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"66",X"00",X"00",X"30",X"60",X"00",X"00",X"30",X"00",X"11",X"00",
		X"00",X"00",X"66",X"33",X"00",X"00",X"01",X"31",X"00",X"00",X"11",X"30",X"00",X"00",X"00",X"3F",
		X"00",X"00",X"11",X"33",X"00",X"00",X"01",X"06",X"00",X"00",X"01",X"06",X"00",X"00",X"10",X"66",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"43",X"33",X"00",X"00",X"33",X"66",X"00",X"00",X"06",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"04",X"01",X"00",X"03",X"34",X"11",X"00",X"00",X"10",X"00",X"00",
		X"06",X"06",X"00",X"00",X"06",X"11",X"60",X"00",X"00",X"01",X"33",X"00",X"00",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"01",X"06",X"11",X"00",X"01",X"00",X"00",X"00",
		X"01",X"01",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"0A",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"0B",X"00",X"0B",X"00",X"AA",X"EE",X"E0",X"00",X"00",X"99",X"F5",
		X"00",X"77",X"F9",X"FF",X"00",X"55",X"9F",X"99",X"00",X"55",X"9F",X"FF",X"00",X"FF",X"9F",X"FF",
		X"00",X"55",X"FF",X"F9",X"00",X"33",X"FF",X"FF",X"B0",X"33",X"FF",X"FF",X"00",X"33",X"FF",X"FF",
		X"0B",X"33",X"FF",X"FF",X"00",X"33",X"FF",X"FF",X"00",X"33",X"FF",X"FF",X"0A",X"55",X"FF",X"F9",
		X"0B",X"FF",X"9F",X"FF",X"0A",X"55",X"9F",X"FF",X"00",X"55",X"9F",X"99",X"00",X"77",X"F9",X"FF",
		X"00",X"00",X"99",X"F5",X"00",X"00",X"EE",X"BB",X"00",X"00",X"AA",X"AA",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"BA",X"00",X"00",X"0B",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"A0",X"0A",X"0B",X"00",X"00",X"A0",X"B0",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"9F",X"99",X"00",X"55",X"9F",X"FF",X"00",X"FF",X"9F",X"FF",
		X"00",X"55",X"FF",X"F9",X"00",X"33",X"FF",X"FF",X"00",X"33",X"FF",X"FF",X"00",X"33",X"FF",X"FF",
		X"00",X"33",X"FF",X"FF",X"00",X"33",X"FF",X"FF",X"00",X"33",X"FF",X"FF",X"00",X"55",X"FF",X"F9",
		X"00",X"FF",X"9F",X"FF",X"00",X"55",X"9F",X"FF",X"00",X"00",X"9F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"A0",X"00",X"0A",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"BB",X"B0",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"A0",X"00",X"BB",X"00",X"0A",X"00",X"B0",X"9F",X"B0",
		X"0B",X"05",X"FF",X"0B",X"00",X"33",X"FF",X"00",X"00",X"53",X"FF",X"00",X"00",X"03",X"FF",X"00",
		X"00",X"00",X"FF",X"0B",X"00",X"33",X"FF",X"0B",X"00",X"00",X"FF",X"0B",X"00",X"05",X"FF",X"00",
		X"00",X"00",X"9F",X"00",X"00",X"55",X"9F",X"0B",X"00",X"00",X"9F",X"0B",X"00",X"B0",X"00",X"BB",
		X"00",X"BB",X"BB",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"0B",X"00",X"B0",X"00",X"B0",X"00",X"0B",
		X"00",X"B0",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"0A",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"0B",
		X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"93",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"B0",X"B0",X"00",X"00",X"B0",X"B0",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"0B",X"00",
		X"BB",X"00",X"0B",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"B0",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"0B",X"0B",X"BB",X"00",X"0B",X"BB",X"BB",X"00",
		X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"B0",X"00",X"0B",X"BB",X"B0",X"0B",X"B0",X"BB",X"B0",X"00",
		X"B0",X"BB",X"00",X"BB",X"BB",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"BB",X"BB",X"B0",X"B0",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"B0",X"B0",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"B0",X"BB",
		X"BB",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"0B",X"00",X"B0",X"BB",X"00",X"BB",
		X"B0",X"BB",X"B0",X"00",X"0B",X"BB",X"B0",X"0B",X"0B",X"BB",X"B0",X"00",X"0B",X"BB",X"BB",X"00",
		X"0B",X"BB",X"BB",X"00",X"0B",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"B0",X"0B",X"BB",X"00",
		X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"0B",X"00",
		X"BB",X"00",X"0B",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"B0",X"B0",X"00",X"00",X"B0",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"49",X"00",
		X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"92",
		X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"99",X"22",X"29",X"22",X"99",X"22",X"29",X"22",X"99",
		X"22",X"29",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",
		X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",
		X"22",X"2A",X"22",X"A9",X"22",X"AA",X"22",X"AA",X"22",X"AA",X"22",X"AA",X"22",X"A9",X"22",X"9A",
		X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"99",X"29",X"92",X"22",X"9E",X"22",X"22",X"22",X"99",X"22",X"22",
		X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"29",X"92",X"22",X"99",X"22",X"22",
		X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"29",X"92",X"22",X"99",X"22",X"22",
		X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"29",X"92",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"29",X"29",X"22",
		X"22",X"92",X"92",X"92",X"22",X"29",X"99",X"22",X"22",X"92",X"99",X"92",X"22",X"29",X"59",X"22",
		X"22",X"92",X"59",X"92",X"22",X"29",X"E5",X"22",X"22",X"92",X"EE",X"92",X"22",X"29",X"FE",X"22",
		X"22",X"92",X"FE",X"92",X"22",X"25",X"EE",X"22",X"22",X"FF",X"E5",X"92",X"22",X"2F",X"5F",X"22",
		X"22",X"92",X"F2",X"92",X"22",X"29",X"29",X"22",X"22",X"92",X"92",X"92",X"22",X"29",X"29",X"22",
		X"22",X"92",X"92",X"92",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"09",X"90",X"90",X"00",
		X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"90",
		X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",
		X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",
		X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",
		X"09",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",
		X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"55",X"00",X"00",X"5F",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"EE",X"00",X"09",X"FE",X"EE",X"00",X"9F",X"EE",X"E9",
		X"00",X"F5",X"EE",X"55",X"00",X"95",X"55",X"99",X"00",X"FF",X"5F",X"9E",X"00",X"FF",X"5F",X"59",
		X"00",X"FF",X"5F",X"55",X"00",X"FF",X"5F",X"55",X"00",X"FE",X"5F",X"55",X"0F",X"FF",X"5F",X"55",
		X"0F",X"FF",X"5F",X"55",X"00",X"EF",X"5F",X"55",X"00",X"FF",X"5F",X"55",X"00",X"55",X"5F",X"55",
		X"00",X"55",X"5F",X"59",X"00",X"FF",X"5F",X"9F",X"00",X"9F",X"5E",X"99",X"00",X"FF",X"E5",X"FF",
		X"00",X"5F",X"55",X"53",X"00",X"05",X"55",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E5",X"99",X"99",X"00",X"55",X"55",X"55",X"00",
		X"FF",X"FF",X"FF",X"00",X"EE",X"FF",X"FF",X"00",X"EE",X"22",X"22",X"00",X"EE",X"42",X"44",X"00",
		X"5F",X"44",X"44",X"00",X"97",X"44",X"44",X"00",X"47",X"44",X"44",X"00",X"47",X"44",X"44",X"00",
		X"47",X"44",X"44",X"00",X"47",X"44",X"44",X"00",X"47",X"44",X"44",X"00",X"44",X"44",X"44",X"00",
		X"24",X"44",X"44",X"00",X"47",X"44",X"44",X"00",X"27",X"44",X"44",X"00",X"42",X"44",X"44",X"00",
		X"27",X"44",X"44",X"00",X"22",X"44",X"44",X"00",X"92",X"24",X"24",X"00",X"F3",X"22",X"22",X"00",
		X"55",X"22",X"22",X"00",X"55",X"FF",X"FF",X"00",X"55",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"E0",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"55",
		X"00",X"99",X"44",X"33",X"00",X"99",X"99",X"99",X"00",X"94",X"99",X"39",X"00",X"49",X"99",X"22",
		X"00",X"99",X"9E",X"22",X"00",X"99",X"E5",X"39",X"09",X"99",X"99",X"93",X"99",X"AA",X"AA",X"33",
		X"09",X"AA",X"FF",X"33",X"00",X"AA",X"AF",X"33",X"00",X"AA",X"AA",X"33",X"00",X"4A",X"AA",X"99",
		X"00",X"A4",X"AA",X"93",X"00",X"AA",X"AA",X"39",X"00",X"9A",X"44",X"99",X"00",X"99",X"AA",X"FF",
		X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"E0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"EE",X"E9",X"00",X"00",
		X"9E",X"E9",X"00",X"00",X"9E",X"E9",X"00",X"00",X"9E",X"E9",X"00",X"00",X"EE",X"39",X"00",X"00",
		X"99",X"99",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",
		X"EE",X"55",X"00",X"00",X"55",X"33",X"00",X"00",X"EE",X"99",X"00",X"00",X"9E",X"E9",X"00",X"00",
		X"9E",X"E9",X"00",X"00",X"9E",X"E9",X"00",X"00",X"EE",X"E9",X"00",X"00",X"5E",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"0C",
		X"00",X"00",X"11",X"00",X"00",X"00",X"99",X"0A",X"00",X"00",X"00",X"F0",X"00",X"90",X"99",X"00",
		X"00",X"40",X"00",X"00",X"00",X"46",X"00",X"0A",X"00",X"40",X"00",X"00",X"00",X"49",X"99",X"00",
		X"00",X"00",X"11",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"CA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"11",X"F0",
		X"00",X"49",X"99",X"00",X"00",X"40",X"00",X"F0",X"00",X"49",X"00",X"E0",X"00",X"40",X"00",X"0A",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"99",X"EB",X"00",X"00",X"11",X"A0",
		X"00",X"00",X"AA",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"50",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"50",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"05",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"50",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"CC",X"CC",X"BC",X"00",X"EB",X"00",X"99",X"00",X"AA",X"BE",X"CC",X"99",X"AC",X"AA",X"BB",
		X"59",X"AA",X"EB",X"0B",X"59",X"BE",X"BE",X"C9",X"4C",X"EB",X"BB",X"BC",X"4C",X"BB",X"B5",X"EB",
		X"0C",X"BB",X"BB",X"BB",X"0C",X"EE",X"5B",X"BB",X"0C",X"5F",X"B5",X"BB",X"0C",X"BB",X"5B",X"BB",
		X"0C",X"BB",X"B5",X"BB",X"4C",X"BB",X"5B",X"BB",X"4C",X"BB",X"BF",X"69",X"50",X"66",X"FB",X"9B",
		X"50",X"BB",X"BB",X"BB",X"00",X"9C",X"6F",X"BB",X"00",X"EB",X"BB",X"CC",X"00",X"BE",X"00",X"99",
		X"00",X"CC",X"CC",X"BC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"97",X"99",X"99",X"00",X"77",X"9D",X"99",
		X"00",X"77",X"DD",X"99",X"00",X"00",X"DD",X"99",X"00",X"99",X"9A",X"E9",X"00",X"91",X"77",X"EE",
		X"9F",X"11",X"D7",X"EE",X"99",X"11",X"7D",X"EE",X"9F",X"1F",X"77",X"EE",X"99",X"1F",X"77",X"EE",
		X"00",X"01",X"77",X"EE",X"00",X"00",X"7D",X"E0",X"00",X"99",X"DD",X"00",X"00",X"77",X"7D",X"00",
		X"00",X"76",X"07",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"A9",X"09",X"5E",X"90",
		X"99",X"99",X"EE",X"90",X"99",X"99",X"99",X"91",X"FF",X"FF",X"F9",X"91",X"99",X"99",X"99",X"44",
		X"9E",X"AA",X"57",X"A1",X"EA",X"AA",X"AA",X"51",X"EA",X"AA",X"AA",X"99",X"AA",X"AA",X"AA",X"AA",
		X"EA",X"94",X"AA",X"AE",X"AA",X"49",X"AA",X"EE",X"EA",X"49",X"AA",X"E5",X"AA",X"A4",X"AA",X"E5",
		X"EA",X"A9",X"AA",X"E5",X"AE",X"94",X"AA",X"E5",X"EA",X"49",X"AA",X"EE",X"EE",X"49",X"AA",X"AE",
		X"EA",X"E4",X"AA",X"AA",X"5E",X"AE",X"AA",X"99",X"E5",X"EE",X"AE",X"51",X"9E",X"EE",X"55",X"A1",
		X"99",X"99",X"99",X"44",X"FF",X"FF",X"F9",X"91",X"99",X"99",X"99",X"91",X"99",X"D9",X"EE",X"99",
		X"D9",X"09",X"0E",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"00",X"00",X"A9",X"31",X"00",X"00",
		X"33",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"55",X"01",X"00",X"00",X"9C",X"10",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"30",X"00",X"00",X"A5",X"90",X"00",X"00",
		X"55",X"A9",X"00",X"00",X"FF",X"A9",X"00",X"00",X"55",X"A9",X"00",X"00",X"55",X"A9",X"00",X"00",
		X"55",X"A9",X"00",X"00",X"A5",X"90",X"00",X"00",X"95",X"30",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"9C",X"10",X"00",X"00",X"55",X"01",X"00",X"00",X"EE",X"11",X"00",X"00",
		X"99",X"41",X"00",X"00",X"A9",X"91",X"00",X"00",X"0E",X"19",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"07",X"01",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"09",X"90",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"AE",X"99",X"99",X"00",X"EE",X"E9",X"99",X"00",X"E5",X"AE",X"AE",
		X"00",X"EE",X"99",X"9A",X"00",X"AA",X"A9",X"A9",X"00",X"99",X"99",X"9A",X"00",X"FF",X"99",X"99",
		X"00",X"FF",X"99",X"7A",X"00",X"99",X"99",X"AE",X"00",X"F9",X"9A",X"EA",X"00",X"F9",X"AA",X"AE",
		X"00",X"F9",X"AE",X"EA",X"00",X"F9",X"AE",X"EE",X"00",X"F9",X"AE",X"EE",X"00",X"F9",X"AE",X"EE",
		X"00",X"F9",X"AA",X"5E",X"00",X"F9",X"9A",X"EE",X"00",X"99",X"99",X"E5",X"00",X"FF",X"99",X"56",
		X"00",X"FF",X"99",X"AA",X"00",X"99",X"99",X"DD",X"00",X"EA",X"99",X"DD",X"00",X"E5",X"E9",X"DD",
		X"00",X"5E",X"EE",X"AA",X"00",X"E5",X"EE",X"EE",X"00",X"EE",X"99",X"09",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"5E",X"99",X"00",X"00",X"99",X"95",X"00",X"00",
		X"9A",X"95",X"00",X"00",X"A9",X"95",X"00",X"00",X"9A",X"95",X"00",X"00",X"99",X"95",X"00",X"00",
		X"7A",X"95",X"00",X"00",X"AA",X"95",X"00",X"00",X"EA",X"95",X"00",X"00",X"AA",X"95",X"00",X"00",
		X"EA",X"95",X"00",X"00",X"AA",X"95",X"00",X"00",X"EA",X"95",X"00",X"00",X"AA",X"95",X"00",X"00",
		X"EA",X"95",X"00",X"00",X"AA",X"95",X"00",X"00",X"EA",X"95",X"00",X"00",X"55",X"95",X"00",X"00",
		X"AA",X"95",X"00",X"00",X"DD",X"95",X"00",X"00",X"DD",X"95",X"00",X"00",X"DD",X"95",X"00",X"00",
		X"AA",X"95",X"00",X"00",X"E5",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"5F",X"FF",X"00",X"11",X"5F",X"55",X"00",X"11",X"5F",X"9A",X"00",X"11",X"5F",X"9A",
		X"00",X"11",X"5F",X"9A",X"00",X"11",X"5F",X"99",X"00",X"22",X"5F",X"F9",X"00",X"92",X"15",X"F9",
		X"00",X"19",X"15",X"F9",X"00",X"12",X"15",X"F9",X"00",X"12",X"15",X"FF",X"00",X"11",X"95",X"F9",
		X"00",X"11",X"15",X"F9",X"00",X"11",X"15",X"FF",X"00",X"11",X"11",X"BF",X"00",X"22",X"21",X"BF",
		X"00",X"11",X"11",X"AF",X"00",X"11",X"99",X"9F",X"00",X"11",X"11",X"9F",X"00",X"11",X"11",X"FF",
		X"00",X"11",X"11",X"55",X"00",X"11",X"11",X"91",X"00",X"12",X"11",X"22",X"00",X"91",X"12",X"12",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"91",X"11",X"11",X"00",X"91",X"11",X"11",
		X"00",X"99",X"91",X"99",X"00",X"00",X"00",X"00",X"00",X"09",X"EE",X"EE",X"00",X"09",X"99",X"99",
		X"00",X"22",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"09",X"22",X"92",X"99",X"90",X"93",X"22",X"22",
		X"02",X"92",X"29",X"22",X"09",X"22",X"22",X"22",X"02",X"22",X"22",X"22",X"02",X"22",X"22",X"22",
		X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"92",X"32",X"33",X"33",X"92",X"39",X"33",X"99",
		X"92",X"33",X"33",X"33",X"92",X"33",X"11",X"33",X"91",X"11",X"11",X"11",X"91",X"11",X"11",X"11",
		X"91",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"11",X"22",X"22",X"01",X"22",X"21",X"11",
		X"09",X"99",X"11",X"11",X"02",X"11",X"11",X"11",X"09",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"11",X"99",X"99",X"00",X"11",X"29",X"29",X"00",X"21",X"99",X"99",X"00",X"11",X"99",X"99",
		X"00",X"39",X"99",X"99",X"00",X"39",X"33",X"EE",X"00",X"33",X"33",X"33",X"00",X"99",X"91",X"99",
		X"00",X"92",X"12",X"22",X"00",X"92",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"92",
		X"00",X"22",X"22",X"99",X"00",X"92",X"22",X"99",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"99",
		X"00",X"22",X"22",X"92",X"00",X"22",X"22",X"92",X"00",X"22",X"22",X"22",X"00",X"12",X"23",X"22",
		X"00",X"29",X"2F",X"22",X"00",X"22",X"2F",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"29",X"99",X"92",X"00",X"22",X"22",X"29",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"29",X"99",X"92",X"00",X"22",X"22",X"29",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",
		X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"22",X"22",X"F3",X"00",X"21",X"22",X"F3",X"00",
		X"21",X"22",X"F3",X"00",X"21",X"91",X"F3",X"00",X"21",X"11",X"F3",X"00",X"91",X"11",X"F3",X"00",
		X"92",X"11",X"F3",X"00",X"92",X"11",X"F3",X"00",X"92",X"22",X"F3",X"00",X"92",X"11",X"F3",X"55",
		X"99",X"11",X"F3",X"55",X"92",X"11",X"F3",X"35",X"92",X"11",X"F3",X"35",X"92",X"21",X"FF",X"35",
		X"92",X"21",X"FF",X"55",X"11",X"21",X"FF",X"55",X"22",X"22",X"FF",X"55",X"11",X"11",X"FF",X"35",
		X"11",X"11",X"9F",X"30",X"11",X"11",X"9F",X"00",X"11",X"11",X"9F",X"00",X"11",X"91",X"9F",X"00",
		X"99",X"99",X"9F",X"00",X"EE",X"EE",X"EE",X"00",X"EE",X"EE",X"9E",X"00",X"EE",X"99",X"9E",X"00",
		X"29",X"99",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",
		X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"92",X"22",X"F3",X"00",X"22",X"99",X"F3",X"00",
		X"22",X"92",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",
		X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"33",X"33",X"F3",X"00",X"99",X"99",X"F3",X"00",
		X"33",X"33",X"F3",X"00",X"11",X"33",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",
		X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"21",X"22",X"F3",X"00",
		X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",
		X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"12",X"F3",X"00",X"22",X"21",X"F3",X"00",
		X"33",X"99",X"93",X"00",X"EE",X"33",X"93",X"00",X"33",X"33",X"33",X"00",X"99",X"99",X"9F",X"00",
		X"11",X"91",X"9F",X"00",X"22",X"22",X"9F",X"00",X"22",X"22",X"9F",X"00",X"22",X"22",X"9F",X"30",
		X"22",X"22",X"FF",X"35",X"99",X"92",X"FF",X"55",X"11",X"12",X"FF",X"55",X"22",X"22",X"FF",X"55",
		X"22",X"22",X"FF",X"35",X"22",X"22",X"F3",X"35",X"22",X"99",X"F3",X"35",X"99",X"22",X"F3",X"55",
		X"22",X"22",X"F3",X"55",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",
		X"92",X"29",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"33",X"F3",X"00",
		X"11",X"32",X"F3",X"00",X"22",X"32",X"F3",X"00",X"29",X"39",X"F3",X"00",X"22",X"92",X"F3",X"00",
		X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",
		X"00",X"00",X"09",X"90",X"00",X"00",X"90",X"99",X"00",X"09",X"99",X"11",X"00",X"00",X"55",X"99",
		X"00",X"99",X"55",X"39",X"00",X"55",X"55",X"39",X"00",X"55",X"55",X"35",X"00",X"55",X"55",X"53",
		X"00",X"55",X"31",X"33",X"00",X"53",X"77",X"77",X"00",X"14",X"33",X"99",X"99",X"47",X"33",X"BB",
		X"00",X"71",X"3A",X"99",X"00",X"55",X"AB",X"99",X"00",X"55",X"AB",X"99",X"00",X"55",X"AB",X"39",
		X"00",X"FF",X"AB",X"59",X"00",X"FF",X"AB",X"99",X"00",X"FF",X"AB",X"99",X"00",X"11",X"5A",X"99",
		X"99",X"41",X"FF",X"BB",X"00",X"11",X"FF",X"FF",X"00",X"55",X"11",X"11",X"00",X"55",X"51",X"55",
		X"00",X"55",X"55",X"55",X"00",X"FF",X"55",X"35",X"00",X"FF",X"55",X"39",X"00",X"00",X"FF",X"39",
		X"00",X"00",X"FF",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"00",X"00",
		X"90",X"99",X"09",X"00",X"99",X"99",X"90",X"00",X"99",X"FF",X"09",X"00",X"59",X"99",X"99",X"00",
		X"55",X"39",X"99",X"00",X"95",X"99",X"90",X"00",X"99",X"F9",X"99",X"00",X"11",X"11",X"39",X"00",
		X"99",X"99",X"F0",X"00",X"99",X"FF",X"09",X"00",X"59",X"99",X"90",X"00",X"59",X"FF",X"09",X"00",
		X"59",X"FF",X"99",X"00",X"59",X"99",X"90",X"00",X"99",X"FF",X"99",X"00",X"99",X"99",X"F0",X"00",
		X"44",X"11",X"00",X"00",X"55",X"FF",X"90",X"00",X"FF",X"99",X"09",X"00",X"FF",X"F9",X"90",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"06",X"00",
		X"90",X"99",X"16",X"00",X"99",X"99",X"66",X"00",X"99",X"F6",X"16",X"60",X"59",X"99",X"96",X"00",
		X"55",X"39",X"99",X"00",X"95",X"99",X"90",X"00",X"99",X"F9",X"99",X"00",X"11",X"11",X"39",X"00",
		X"99",X"99",X"F0",X"00",X"99",X"FF",X"09",X"00",X"59",X"99",X"90",X"00",X"59",X"FF",X"09",X"00",
		X"59",X"FF",X"99",X"00",X"59",X"99",X"90",X"00",X"99",X"FF",X"99",X"00",X"99",X"99",X"F0",X"00",
		X"44",X"11",X"00",X"00",X"55",X"FF",X"90",X"00",X"FF",X"99",X"09",X"00",X"FF",X"F9",X"90",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"99",X"60",X"F0",X"00",X"90",X"66",X"00",X"00",X"F6",X"FF",X"00",
		X"00",X"01",X"61",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"00",X"00",
		X"90",X"99",X"09",X"00",X"99",X"99",X"90",X"60",X"99",X"FF",X"06",X"00",X"59",X"99",X"99",X"00",
		X"55",X"39",X"99",X"00",X"95",X"99",X"90",X"00",X"99",X"F9",X"99",X"00",X"11",X"11",X"39",X"00",
		X"99",X"99",X"F0",X"00",X"99",X"FF",X"09",X"00",X"59",X"99",X"90",X"00",X"59",X"FF",X"09",X"00",
		X"59",X"FF",X"99",X"00",X"59",X"99",X"90",X"00",X"99",X"FF",X"99",X"00",X"99",X"99",X"F0",X"00",
		X"44",X"11",X"00",X"00",X"55",X"FF",X"90",X"00",X"FF",X"99",X"09",X"00",X"FF",X"F9",X"90",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"99",X"06",X"00",X"00",X"90",X"66",X"00",X"00",X"F0",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"22",X"90",X"00",X"00",X"AA",X"10",X"00",X"00",X"11",X"90",X"00",X"00",
		X"11",X"10",X"00",X"00",X"11",X"90",X"00",X"00",X"92",X"10",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"10",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"90",X"00",X"00",
		X"99",X"10",X"00",X"00",X"99",X"90",X"00",X"00",X"92",X"10",X"00",X"00",X"11",X"90",X"00",X"00",
		X"11",X"10",X"00",X"00",X"1F",X"00",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"5E",X"99",X"00",X"00",X"99",X"95",X"00",X"00",
		X"9A",X"95",X"00",X"00",X"A9",X"95",X"00",X"00",X"9A",X"91",X"00",X"00",X"99",X"15",X"00",X"00",
		X"7A",X"11",X"00",X"00",X"AA",X"15",X"00",X"00",X"EA",X"91",X"00",X"00",X"AA",X"95",X"00",X"00",
		X"EA",X"95",X"00",X"00",X"AA",X"95",X"00",X"00",X"EA",X"95",X"00",X"00",X"AA",X"95",X"00",X"00",
		X"EA",X"95",X"00",X"00",X"AA",X"91",X"00",X"00",X"EA",X"15",X"00",X"00",X"55",X"11",X"00",X"00",
		X"AA",X"15",X"00",X"00",X"DD",X"91",X"00",X"00",X"DD",X"95",X"00",X"00",X"DD",X"95",X"00",X"00",
		X"AA",X"95",X"00",X"00",X"E5",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"92",X"22",X"00",X"00",X"21",X"11",
		X"00",X"00",X"11",X"10",X"00",X"00",X"77",X"22",X"00",X"00",X"29",X"29",X"00",X"01",X"92",X"92",
		X"00",X"11",X"99",X"99",X"00",X"17",X"44",X"44",X"00",X"72",X"44",X"44",X"00",X"22",X"44",X"94",
		X"00",X"22",X"44",X"49",X"00",X"22",X"46",X"94",X"00",X"22",X"66",X"29",X"0C",X"22",X"69",X"22",
		X"CC",X"22",X"99",X"22",X"C6",X"92",X"99",X"22",X"CC",X"29",X"99",X"24",X"0C",X"92",X"69",X"44",
		X"06",X"29",X"F3",X"44",X"00",X"92",X"7F",X"44",X"00",X"99",X"77",X"44",X"00",X"29",X"44",X"44",
		X"00",X"29",X"46",X"44",X"00",X"11",X"22",X"92",X"00",X"11",X"99",X"29",X"00",X"67",X"92",X"92",
		X"00",X"01",X"29",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"11",X"11",X"00",X"00",X"77",X"72",
		X"00",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"22",X"99",X"09",X"00",X"10",X"22",X"99",X"00",
		X"11",X"11",X"22",X"00",X"12",X"11",X"11",X"00",X"22",X"21",X"11",X"90",X"92",X"92",X"92",X"09",
		X"22",X"99",X"29",X"90",X"22",X"79",X"92",X"99",X"22",X"79",X"99",X"29",X"22",X"79",X"62",X"29",
		X"22",X"79",X"29",X"29",X"22",X"79",X"62",X"19",X"22",X"72",X"29",X"29",X"22",X"22",X"62",X"19",
		X"22",X"22",X"29",X"29",X"22",X"22",X"62",X"19",X"22",X"22",X"29",X"29",X"22",X"22",X"62",X"10",
		X"22",X"22",X"29",X"20",X"22",X"22",X"62",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"29",X"00",
		X"22",X"22",X"92",X"00",X"22",X"29",X"29",X"00",X"29",X"99",X"21",X"00",X"99",X"92",X"11",X"00",
		X"21",X"11",X"12",X"00",X"11",X"11",X"00",X"00",X"11",X"20",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"05",X"00",X"00",X"F0",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"50",X"F5",X"00",
		X"55",X"50",X"55",X"00",X"55",X"05",X"55",X"00",X"00",X"55",X"50",X"00",X"00",X"50",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"50",X"00",X"5F",X"F5",X"55",
		X"55",X"55",X"05",X"F0",X"00",X"55",X"50",X"FF",X"00",X"55",X"00",X"05",X"00",X"05",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"50",X"05",X"00",X"00",X"05",X"55",X"00",X"00",X"50",X"55",X"00",
		X"00",X"5F",X"50",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"05",X"55",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",
		X"00",X"0F",X"05",X"00",X"00",X"F0",X"55",X"00",X"00",X"55",X"50",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"F5",X"05",X"00",X"00",X"5F",X"50",X"00",X"00",X"05",X"05",X"00",
		X"00",X"00",X"55",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",
		X"90",X"15",X"50",X"00",X"99",X"F1",X"55",X"00",X"99",X"11",X"55",X"00",X"F9",X"11",X"55",X"00",
		X"F9",X"11",X"55",X"00",X"F5",X"55",X"55",X"00",X"FF",X"55",X"55",X"00",X"FF",X"55",X"55",X"00",
		X"FF",X"F5",X"15",X"50",X"FF",X"FF",X"11",X"55",X"0F",X"F3",X"11",X"55",X"0F",X"F3",X"11",X"55",
		X"0F",X"F3",X"31",X"11",X"0F",X"F3",X"5F",X"11",X"0F",X"F3",X"9F",X"19",X"00",X"FF",X"BB",X"99",
		X"00",X"1F",X"9B",X"99",X"00",X"1F",X"99",X"59",X"00",X"11",X"99",X"55",X"00",X"11",X"91",X"25",
		X"00",X"11",X"51",X"25",X"00",X"11",X"51",X"25",X"00",X"51",X"55",X"22",X"00",X"51",X"95",X"22",
		X"00",X"51",X"99",X"12",X"00",X"51",X"B9",X"91",X"00",X"51",X"BB",X"33",X"00",X"51",X"FB",X"F3",
		X"55",X"11",X"5F",X"99",X"05",X"51",X"FF",X"99",X"05",X"55",X"FF",X"FF",X"00",X"F5",X"3F",X"F0",
		X"00",X"0F",X"9F",X"FF",X"00",X"00",X"99",X"19",X"00",X"99",X"19",X"99",X"00",X"09",X"11",X"3F",
		X"00",X"00",X"F1",X"31",X"00",X"00",X"F1",X"99",X"00",X"00",X"9F",X"F9",X"00",X"00",X"90",X"FF",
		X"00",X"00",X"90",X"FF",X"00",X"00",X"90",X"FF",X"00",X"00",X"90",X"FF",X"00",X"00",X"90",X"FF",
		X"00",X"00",X"99",X"3F",X"00",X"00",X"99",X"39",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"09",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"99",X"99",X"DD",X"00",X"00",X"09",X"BB",X"00",X"00",X"09",X"99",
		X"00",X"00",X"99",X"00",X"00",X"09",X"DD",X"00",X"00",X"9B",X"99",X"00",X"00",X"BF",X"B9",X"00",
		X"00",X"4B",X"99",X"90",X"90",X"4F",X"BB",X"99",X"00",X"4B",X"BB",X"B9",X"00",X"49",X"FB",X"BB",
		X"00",X"44",X"BF",X"BB",X"00",X"4F",X"FB",X"BB",X"00",X"4F",X"BF",X"BB",X"F0",X"4F",X"FB",X"BB",
		X"00",X"4F",X"BF",X"BB",X"00",X"49",X"FB",X"BB",X"00",X"44",X"BF",X"BB",X"00",X"4B",X"FB",X"FB",
		X"00",X"4F",X"BF",X"BA",X"90",X"4F",X"FB",X"99",X"00",X"4F",X"B9",X"90",X"00",X"FF",X"B9",X"00",
		X"00",X"AF",X"99",X"00",X"00",X"0B",X"AA",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"09",X"99",
		X"00",X"00",X"09",X"DD",X"00",X"99",X"99",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"B0",X"00",X"00",X"0A",X"B9",X"A9",X"00",X"0A",
		X"B9",X"DB",X"9A",X"09",X"B9",X"BD",X"BD",X"99",X"B9",X"BB",X"BB",X"BB",X"B9",X"FF",X"FF",X"BB",
		X"59",X"55",X"B5",X"BB",X"B9",X"BB",X"BB",X"AB",X"B9",X"DB",X"AA",X"0F",X"B9",X"AA",X"00",X"0B",
		X"B0",X"00",X"00",X"0B",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"AA",X"00",X"00",X"22",X"49",X"00",X"00",X"22",X"49",X"00",X"00",X"22",X"49",X"00",
		X"00",X"2B",X"F9",X"DD",X"00",X"BB",X"F4",X"0D",X"00",X"BB",X"F4",X"0B",X"00",X"BB",X"B9",X"00",
		X"00",X"FF",X"44",X"00",X"00",X"9B",X"FF",X"90",X"00",X"AF",X"FF",X"D9",X"00",X"B9",X"F4",X"D9",
		X"00",X"B4",X"94",X"D9",X"00",X"4F",X"4F",X"99",X"00",X"FF",X"4B",X"99",X"00",X"FF",X"FF",X"BA",
		X"00",X"BF",X"FB",X"BA",X"00",X"B4",X"BF",X"B9",X"00",X"9B",X"FB",X"99",X"00",X"99",X"9F",X"99",
		X"00",X"00",X"A9",X"99",X"00",X"00",X"AA",X"9A",X"00",X"90",X"AA",X"9B",X"00",X"99",X"0A",X"9B",
		X"00",X"09",X"00",X"9B",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"BB",X"9E",
		X"00",X"00",X"BB",X"0E",X"00",X"00",X"BB",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"BD",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"D0",X"00",X"00",X"BB",X"BD",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"DB",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"BF",X"00",X"D0",X"00",X"BB",X"D0",X"DD",X"00",X"DB",X"BD",X"DD",X"00",X"0D",X"BB",X"BB",
		X"00",X"00",X"FB",X"AB",X"00",X"00",X"FF",X"AA",X"00",X"00",X"BF",X"AA",X"00",X"00",X"DB",X"AA",
		X"00",X"00",X"0D",X"A0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"02",X"94",X"00",X"00",
		X"22",X"94",X"09",X"00",X"22",X"4D",X"09",X"00",X"22",X"4F",X"99",X"00",X"BB",X"49",X"00",X"00",
		X"BB",X"A9",X"00",X"00",X"BB",X"49",X"90",X"00",X"BB",X"44",X"D9",X"00",X"B4",X"FF",X"99",X"00",
		X"A4",X"FF",X"D9",X"00",X"49",X"FF",X"D9",X"00",X"AB",X"9F",X"DD",X"00",X"A4",X"F9",X"9D",X"00",
		X"44",X"94",X"DD",X"00",X"A4",X"44",X"9D",X"0D",X"AB",X"5F",X"9D",X"D9",X"AB",X"FB",X"9D",X"D9",
		X"AA",X"BF",X"99",X"D9",X"0A",X"FB",X"A9",X"DD",X"0A",X"BF",X"B9",X"BD",X"99",X"FB",X"99",X"BB",
		X"99",X"9F",X"B9",X"9B",X"90",X"9B",X"99",X"9B",X"90",X"99",X"9B",X"90",X"99",X"99",X"BB",X"00",
		X"99",X"99",X"B9",X"00",X"09",X"99",X"F9",X"00",X"00",X"0B",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"BA",X"00",X"00",X"00",X"9A",X"00",X"00",X"09",X"AB",X"00",X"00",X"99",X"AB",X"00",
		X"00",X"99",X"AB",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"0A",X"00",X"00",X"99",X"0D",X"00",
		X"00",X"D0",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"D9",X"00",X"D0",X"00",X"DD",X"00",X"D0",
		X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"5B",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",
		X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FB",X"00",
		X"00",X"00",X"FD",X"00",X"00",X"00",X"FD",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"FD",X"00",
		X"00",X"A0",X"B9",X"0D",X"00",X"A0",X"BD",X"0D",X"00",X"AB",X"B9",X"BD",X"00",X"AB",X"FD",X"BD",
		X"00",X"AB",X"F9",X"BD",X"00",X"A0",X"FA",X"0D",X"00",X"00",X"F9",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"0A",X"99",X"00",X"00",X"0A",X"BB",X"00",X"00",X"AA",X"BB",X"90",X"00",X"9A",X"BB",X"90",
		X"00",X"94",X"44",X"99",X"00",X"9F",X"FF",X"90",X"00",X"99",X"FF",X"90",X"00",X"94",X"FF",X"90",
		X"00",X"9A",X"FF",X"90",X"00",X"9A",X"FF",X"90",X"00",X"AA",X"99",X"90",X"00",X"9A",X"44",X"90",
		X"00",X"AA",X"FB",X"90",X"00",X"9A",X"BF",X"99",X"00",X"9A",X"FB",X"90",X"00",X"AA",X"BB",X"90",
		X"00",X"0A",X"BB",X"00",X"00",X"09",X"BB",X"00",X"00",X"09",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",
		X"00",X"99",X"BB",X"99",X"00",X"99",X"F9",X"99",X"00",X"99",X"F9",X"99",X"00",X"99",X"F9",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"A9",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"04",X"00",X"00",X"66",X"06",
		X"00",X"00",X"06",X"60",X"00",X"06",X"00",X"00",X"00",X"06",X"40",X"40",X"00",X"00",X"66",X"60",
		X"00",X"00",X"60",X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"04",X"00",X"46",X"66",X"60",
		X"00",X"66",X"64",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"06",X"00",X"00",X"04",X"60",
		X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"40",X"46",X"00",
		X"00",X"64",X"04",X"40",X"00",X"06",X"00",X"04",X"00",X"00",X"06",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"64",X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"04",X"64",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"64",X"66",X"46",X"00",X"66",X"06",X"66",
		X"00",X"66",X"00",X"60",X"00",X"66",X"00",X"00",X"00",X"06",X"40",X"40",X"00",X"00",X"00",X"60",
		X"04",X"00",X"00",X"04",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"66",X"60",
		X"00",X"00",X"64",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"66",X"04",X"00",X"00",X"04",X"60",
		X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"04",X"66",X"00",X"00",X"46",X"46",X"66",
		X"00",X"66",X"04",X"66",X"00",X"66",X"00",X"06",X"00",X"00",X"06",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"64",X"06",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"00",X"04",X"40",X"00",X"00",X"66",X"64",X"00",X"00",X"60",X"66",X"00",
		X"00",X"44",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"46",X"00",X"66",X"46",X"64",
		X"00",X"66",X"66",X"60",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"40",X"06",X"00",X"04",X"60",
		X"06",X"00",X"00",X"04",X"00",X"00",X"40",X"00",X"00",X"66",X"64",X"04",X"00",X"06",X"66",X"60",
		X"00",X"06",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"66",X"04",X"04",X"00",X"66",X"60",
		X"06",X"00",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"64",X"66",X"00",X"00",X"66",X"46",X"66",
		X"00",X"66",X"04",X"64",X"00",X"66",X"00",X"04",X"00",X"00",X"66",X"00",X"00",X"44",X"04",X"60",
		X"00",X"66",X"04",X"06",X"00",X"06",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"40",X"00",X"40",X"00",X"66",X"00",X"00",X"00",X"60",X"00",X"00",X"04",X"00",X"00",X"00",
		X"00",X"44",X"00",X"04",X"06",X"40",X"00",X"46",X"00",X"60",X"00",X"66",X"00",X"40",X"46",X"66",
		X"00",X"06",X"66",X"60",X"00",X"00",X"66",X"00",X"04",X"00",X"60",X"40",X"66",X"00",X"04",X"66",
		X"06",X"00",X"00",X"66",X"00",X"40",X"40",X"60",X"00",X"66",X"00",X"04",X"00",X"66",X"66",X"60",
		X"00",X"66",X"66",X"00",X"00",X"60",X"06",X"00",X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"66",
		X"06",X"00",X"46",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"40",X"46",X"66",
		X"00",X"64",X"04",X"66",X"00",X"60",X"00",X"06",X"00",X"00",X"00",X"40",X"06",X"44",X"04",X"60",
		X"00",X"66",X"04",X"66",X"00",X"66",X"40",X"66",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"0A",
		X"00",X"0A",X"A0",X"AF",X"00",X"A0",X"0A",X"00",X"00",X"0A",X"A0",X"F0",X"00",X"A0",X"0F",X"00",
		X"0A",X"FA",X"F0",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",X"0A",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"0A",X"00",X"00",X"00",X"A0",X"0A",X"00",X"00",X"0A",X"A0",X"00",
		X"00",X"00",X"0A",X"00",X"0F",X"0A",X"A0",X"A0",X"00",X"F0",X"00",X"00",X"00",X"0F",X"0F",X"A0",
		X"00",X"00",X"F0",X"0A",X"00",X"00",X"00",X"A0",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"0A",X"A0",X"0A",
		X"00",X"A0",X"0A",X"F0",X"00",X"0A",X"AF",X"0F",X"00",X"0F",X"00",X"00",X"0A",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"A0",X"0F",X"0A",X"00",X"00",X"00",X"A0",X"0A",X"00",X"00",X"0A",X"A0",X"00",
		X"00",X"F0",X"0A",X"00",X"00",X"00",X"F0",X"A0",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"FF",X"00",X"F0",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"0F",X"FF",X"F0",X"00",X"FF",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"00",X"F0",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"FF",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"FF",X"00",X"F0",X"FF",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"F0",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"39",X"39",X"93",X"00",X"B3",X"B3",X"3B",X"00",X"B5",X"5B",X"BB",
		X"00",X"FB",X"5F",X"5F",X"00",X"B3",X"B3",X"3B",X"00",X"39",X"39",X"93",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"39",X"39",X"93",X"00",X"B3",X"B3",X"35",X"00",X"B5",X"55",X"55",
		X"00",X"FB",X"5F",X"5F",X"00",X"B3",X"B3",X"35",X"00",X"39",X"39",X"93",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"93",X"00",X"00",X"09",X"30",X"90",X"05",X"90",X"05",X"03",X"50",
		X"95",X"05",X"00",X"00",X"00",X"30",X"30",X"F0",X"00",X"03",X"00",X"00",X"50",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"93",X"00",X"00",X"09",X"30",X"90",X"00",X"90",X"05",X"03",X"00",
		X"95",X"05",X"00",X"F0",X"00",X"30",X"30",X"00",X"00",X"03",X"00",X"50",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"99",X"99",
		X"00",X"09",X"DD",X"99",X"00",X"99",X"D9",X"99",X"00",X"DD",X"99",X"EE",X"00",X"99",X"EE",X"99",
		X"00",X"DD",X"9E",X"55",X"00",X"99",X"9E",X"99",X"00",X"DD",X"9E",X"9E",X"00",X"99",X"EE",X"59",
		X"00",X"DD",X"E5",X"55",X"09",X"99",X"EB",X"55",X"00",X"DD",X"E5",X"55",X"09",X"99",X"EB",X"55",
		X"0A",X"AA",X"B5",X"55",X"0A",X"AB",X"BB",X"55",X"00",X"BA",X"B5",X"55",X"00",X"AB",X"BB",X"55",
		X"00",X"BA",X"BB",X"59",X"00",X"AB",X"A5",X"9F",X"00",X"BA",X"9B",X"99",X"00",X"AB",X"9B",X"55",
		X"00",X"BA",X"B5",X"59",X"00",X"AB",X"55",X"55",X"00",X"BA",X"BA",X"AA",X"00",X"0B",X"AB",X"BB",
		X"00",X"00",X"BA",X"AA",X"00",X"00",X"AB",X"BB",X"00",X"00",X"BA",X"BA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"9D",X"9D",X"00",
		X"99",X"DD",X"9D",X"00",X"99",X"9D",X"99",X"00",X"EE",X"BB",X"55",X"00",X"99",X"DD",X"DD",X"00",
		X"59",X"BB",X"BB",X"00",X"9E",X"DD",X"DD",X"00",X"59",X"BB",X"BB",X"00",X"EA",X"DD",X"DD",X"00",
		X"59",X"BB",X"BB",X"00",X"EA",X"DB",X"DB",X"00",X"E9",X"BB",X"BB",X"00",X"59",X"BB",X"BB",X"00",
		X"EA",X"BA",X"BB",X"00",X"59",X"BB",X"BB",X"00",X"E9",X"AB",X"AB",X"00",X"E9",X"BB",X"BB",X"00",
		X"59",X"AA",X"AA",X"00",X"59",X"BB",X"BB",X"00",X"59",X"AA",X"AA",X"00",X"55",X"BB",X"BB",X"00",
		X"55",X"AA",X"55",X"00",X"55",X"BB",X"9B",X"00",X"AA",X"AA",X"AA",X"00",X"BB",X"BA",X"AA",X"00",
		X"AA",X"AA",X"AA",X"00",X"AB",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"9A",X"9A",X"00",X"0B",X"AB",X"9B",X"00",X"05",X"BD",X"9D",X"00",X"0F",X"BB",X"9B",
		X"00",X"05",X"5B",X"5B",X"00",X"05",X"BA",X"9A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"0A",X"BA",X"9A",
		X"00",X"0B",X"AB",X"AB",X"00",X"05",X"BB",X"9B",X"00",X"0F",X"B5",X"95",X"00",X"05",X"AB",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"F0",X"00",X"FF",X"0F",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"00",
		X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"05",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"FF",X"00",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"F0",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"F0",X"00",X"F0",X"F0",X"0F",
		X"00",X"00",X"0F",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"F0",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"0F",X"0F",X"00",X"F0",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"05",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"05",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"99",X"FA",X"00",X"00",X"59",X"10",X"00",X"00",X"99",X"11",
		X"00",X"09",X"55",X"11",X"00",X"99",X"55",X"11",X"00",X"99",X"55",X"19",X"00",X"99",X"33",X"19",
		X"00",X"09",X"44",X"77",X"00",X"19",X"39",X"93",X"00",X"44",X"33",X"BB",X"00",X"55",X"33",X"99",
		X"00",X"F1",X"35",X"99",X"00",X"11",X"55",X"99",X"00",X"99",X"55",X"99",X"00",X"99",X"55",X"99",
		X"00",X"11",X"59",X"11",X"00",X"31",X"39",X"11",X"00",X"95",X"99",X"11",X"00",X"49",X"99",X"15",
		X"00",X"19",X"19",X"55",X"00",X"99",X"44",X"99",X"00",X"99",X"55",X"19",X"00",X"9F",X"55",X"19",
		X"00",X"9F",X"55",X"19",X"00",X"90",X"F5",X"19",X"00",X"00",X"99",X"19",X"00",X"00",X"F9",X"11",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"F0",X"00",
		X"99",X"99",X"0F",X"00",X"55",X"9F",X"0F",X"F0",X"35",X"FE",X"00",X"0F",X"33",X"33",X"F3",X"0F",
		X"33",X"55",X"33",X"00",X"43",X"93",X"33",X"0F",X"54",X"33",X"33",X"00",X"99",X"33",X"03",X"F0",
		X"F5",X"33",X"30",X"F0",X"55",X"36",X"00",X"00",X"55",X"66",X"00",X"F0",X"55",X"9F",X"00",X"F0",
		X"55",X"9F",X"00",X"0F",X"5F",X"FF",X"00",X"F0",X"99",X"99",X"00",X"0F",X"11",X"41",X"00",X"00",
		X"4F",X"5F",X"00",X"0F",X"FF",X"FF",X"00",X"00",X"55",X"E0",X"00",X"00",X"55",X"9E",X"0F",X"00",
		X"FF",X"99",X"0F",X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"51",
		X"00",X"00",X"55",X"00",X"00",X"99",X"59",X"11",X"00",X"99",X"55",X"11",X"00",X"99",X"53",X"11",
		X"00",X"09",X"34",X"77",X"00",X"99",X"43",X"99",X"00",X"99",X"93",X"BB",X"00",X"59",X"33",X"99",
		X"00",X"FF",X"33",X"99",X"00",X"81",X"35",X"99",X"00",X"19",X"55",X"99",X"00",X"91",X"55",X"99",
		X"00",X"91",X"39",X"99",X"00",X"93",X"99",X"99",X"00",X"95",X"99",X"99",X"00",X"94",X"99",X"91",
		X"00",X"99",X"91",X"11",X"00",X"99",X"54",X"11",X"00",X"99",X"55",X"55",X"00",X"09",X"55",X"15",
		X"00",X"09",X"55",X"99",X"00",X"09",X"99",X"11",X"00",X"00",X"99",X"51",X"00",X"00",X"89",X"F1",
		X"00",X"00",X"09",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"0F",X"00",X"F0",X"F0",X"00",X"0F",X"F0",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"55",X"90",X"00",X"0F",X"33",X"00",X"F0",X"00",X"33",X"0F",X"00",X"00",
		X"73",X"00",X"33",X"F0",X"34",X"0F",X"33",X"00",X"35",X"00",X"33",X"00",X"99",X"30",X"30",X"0F",
		X"9F",X"30",X"03",X"0F",X"95",X"33",X"00",X"00",X"95",X"F6",X"00",X"0F",X"95",X"F9",X"00",X"0F",
		X"95",X"F9",X"00",X"00",X"95",X"FF",X"00",X"0F",X"99",X"99",X"00",X"00",X"31",X"14",X"00",X"00",
		X"54",X"55",X"00",X"00",X"1F",X"9F",X"00",X"F0",X"55",X"9E",X"00",X"00",X"55",X"99",X"00",X"F0",
		X"FF",X"F9",X"00",X"00",X"00",X"0F",X"00",X"F0",X"0F",X"F0",X"00",X"0F",X"00",X"0F",X"FF",X"F0",
		X"0F",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"0F",X"00",X"00",X"00",X"F0",X"55",X"10",X"00",X"00",X"55",X"11",
		X"00",X"99",X"53",X"11",X"00",X"00",X"34",X"77",X"00",X"91",X"43",X"99",X"00",X"99",X"93",X"BB",
		X"00",X"55",X"33",X"90",X"00",X"FF",X"33",X"00",X"0F",X"89",X"35",X"00",X"00",X"19",X"55",X"00",
		X"00",X"99",X"55",X"99",X"00",X"91",X"35",X"99",X"00",X"93",X"39",X"99",X"00",X"95",X"F9",X"99",
		X"00",X"94",X"F9",X"99",X"00",X"99",X"11",X"FF",X"00",X"99",X"54",X"51",X"00",X"99",X"95",X"5F",
		X"00",X"09",X"55",X"55",X"00",X"09",X"99",X"55",X"00",X"09",X"99",X"11",X"00",X"00",X"99",X"51",
		X"00",X"00",X"89",X"F1",X"00",X"00",X"09",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",
		X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",
		X"0F",X"00",X"00",X"00",X"70",X"00",X"00",X"F0",X"30",X"0F",X"00",X"00",X"30",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"F0",X"00",X"00",
		X"95",X"FF",X"00",X"00",X"95",X"0F",X"00",X"00",X"95",X"F0",X"00",X"00",X"99",X"FF",X"00",X"00",
		X"31",X"FF",X"00",X"00",X"54",X"00",X"00",X"00",X"1F",X"FF",X"00",X"F0",X"55",X"00",X"00",X"00",
		X"55",X"0F",X"00",X"F0",X"9F",X"F0",X"00",X"00",X"90",X"00",X"00",X"F0",X"0F",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"0F",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"09",X"55",X"00",X"00",X"55",X"51",
		X"00",X"00",X"55",X"11",X"00",X"F0",X"33",X"77",X"0F",X"00",X"44",X"33",X"00",X"00",X"73",X"AB",
		X"00",X"00",X"33",X"BB",X"00",X"00",X"55",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"33",X"00",
		X"0F",X"00",X"53",X"00",X"0F",X"00",X"F3",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"99",
		X"00",X"00",X"1F",X"99",X"0F",X"00",X"00",X"FF",X"0F",X"00",X"00",X"55",X"0F",X"00",X"00",X"55",
		X"00",X"00",X"09",X"55",X"00",X"0F",X"09",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",
		X"0D",X"F0",X"00",X"00",X"0D",X"FF",X"00",X"00",X"0D",X"00",X"00",X"00",X"DD",X"0F",X"00",X"00",
		X"DD",X"F0",X"00",X"00",X"DD",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"99",X"99",X"F0",X"00",
		X"39",X"99",X"F0",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"09",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"90",X"00",X"00",X"55",X"39",X"09",X"00",X"55",X"33",X"90",X"99",X"15",X"FF",X"00",
		X"00",X"11",X"F5",X"00",X"09",X"11",X"55",X"90",X"09",X"51",X"55",X"90",X"09",X"5F",X"55",X"99",
		X"99",X"55",X"15",X"99",X"99",X"55",X"99",X"11",X"09",X"59",X"99",X"19",X"09",X"59",X"99",X"99",
		X"09",X"F9",X"99",X"99",X"00",X"F9",X"B9",X"95",X"05",X"FF",X"99",X"5F",X"09",X"FF",X"99",X"15",
		X"09",X"1F",X"99",X"11",X"09",X"91",X"99",X"91",X"09",X"91",X"99",X"99",X"00",X"91",X"B9",X"DF",
		X"00",X"95",X"9B",X"DF",X"00",X"5F",X"1F",X"FF",X"00",X"55",X"11",X"FF",X"00",X"5F",X"11",X"F9",
		X"00",X"5F",X"19",X"99",X"00",X"FF",X"19",X"19",X"00",X"FF",X"19",X"F9",X"00",X"FF",X"19",X"F9",
		X"00",X"99",X"19",X"F9",X"00",X"00",X"19",X"FF",X"00",X"00",X"19",X"FF",X"00",X"00",X"19",X"0F",
		X"00",X"11",X"00",X"00",X"09",X"11",X"00",X"00",X"09",X"1F",X"00",X"90",X"00",X"F9",X"00",X"90",
		X"00",X"99",X"19",X"F0",X"00",X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"9F",X"00",
		X"00",X"00",X"FF",X"90",X"00",X"99",X"00",X"90",X"00",X"FF",X"E0",X"F0",X"00",X"99",X"33",X"00",
		X"00",X"99",X"55",X"30",X"00",X"9F",X"59",X"95",X"00",X"11",X"11",X"11",X"00",X"91",X"11",X"99",
		X"00",X"09",X"FF",X"FF",X"00",X"99",X"F9",X"00",X"00",X"F9",X"F9",X"00",X"00",X"FF",X"F9",X"00",
		X"00",X"FF",X"F9",X"00",X"00",X"F9",X"FF",X"FF",X"00",X"9F",X"99",X"99",X"00",X"99",X"11",X"11",
		X"00",X"91",X"11",X"50",X"00",X"99",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"90",
		X"00",X"00",X"99",X"90",X"00",X"FF",X"99",X"F0",X"00",X"9F",X"FF",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"CC",X"99",X"99",
		X"00",X"92",X"22",X"99",X"00",X"29",X"22",X"22",X"00",X"92",X"2C",X"22",X"00",X"99",X"99",X"99",
		X"09",X"29",X"29",X"22",X"09",X"99",X"92",X"22",X"09",X"22",X"92",X"22",X"09",X"22",X"99",X"99",
		X"09",X"C2",X"2C",X"99",X"09",X"22",X"C2",X"92",X"09",X"92",X"22",X"22",X"00",X"99",X"29",X"29",
		X"00",X"C2",X"99",X"99",X"00",X"22",X"22",X"92",X"00",X"C2",X"22",X"22",X"00",X"22",X"22",X"C2",
		X"00",X"99",X"99",X"22",X"00",X"CC",X"22",X"9C",X"00",X"CC",X"2C",X"C9",X"00",X"CC",X"22",X"22",
		X"00",X"22",X"22",X"22",X"09",X"99",X"2C",X"29",X"00",X"C9",X"99",X"99",X"00",X"CC",X"22",X"99",
		X"00",X"22",X"2C",X"99",X"00",X"2C",X"22",X"C9",X"00",X"22",X"22",X"C9",X"00",X"22",X"22",X"C9",
		X"99",X"99",X"99",X"FF",X"22",X"22",X"22",X"F0",X"22",X"22",X"22",X"00",X"99",X"99",X"99",X"00",
		X"22",X"22",X"22",X"90",X"22",X"22",X"22",X"92",X"22",X"22",X"29",X"92",X"99",X"99",X"99",X"29",
		X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"29",X"92",X"99",X"99",X"99",X"F0",
		X"99",X"00",X"F0",X"FF",X"99",X"99",X"F0",X"00",X"22",X"92",X"0F",X"F0",X"2C",X"29",X"02",X"00",
		X"22",X"22",X"20",X"00",X"9C",X"99",X"02",X"00",X"22",X"22",X"90",X"00",X"92",X"29",X"22",X"00",
		X"22",X"92",X"20",X"00",X"99",X"99",X"02",X"00",X"29",X"99",X"20",X"00",X"C2",X"22",X"02",X"00",
		X"92",X"C2",X"20",X"00",X"22",X"9C",X"22",X"F0",X"99",X"22",X"20",X"00",X"99",X"C9",X"02",X"00",
		X"33",X"22",X"20",X"00",X"33",X"22",X"02",X"00",X"39",X"92",X"20",X"00",X"33",X"22",X"02",X"00",
		X"00",X"C9",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"C2",X"22",X"22",
		X"00",X"C2",X"22",X"22",X"00",X"99",X"99",X"99",X"00",X"22",X"99",X"92",X"00",X"22",X"90",X"92",
		X"00",X"22",X"09",X"92",X"00",X"C2",X"90",X"22",X"00",X"C9",X"99",X"99",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"92",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"C2",X"22",X"33",
		X"00",X"C9",X"99",X"29",X"00",X"3C",X"22",X"22",X"00",X"39",X"CC",X"22",X"00",X"39",X"92",X"92",
		X"00",X"39",X"29",X"99",X"00",X"39",X"99",X"00",X"00",X"99",X"F0",X"00",X"0F",X"99",X"2F",X"00",
		X"0F",X"92",X"00",X"00",X"00",X"29",X"02",X"00",X"00",X"99",X"2F",X"00",X"00",X"00",X"F2",X"00",
		X"00",X"0F",X"02",X"00",X"00",X"00",X"2F",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",
		X"99",X"99",X"02",X"00",X"92",X"29",X"20",X"00",X"22",X"92",X"02",X"00",X"29",X"22",X"20",X"00",
		X"C2",X"92",X"22",X"00",X"C9",X"39",X"00",X"F0",X"92",X"92",X"22",X"00",X"22",X"22",X"20",X"00",
		X"92",X"29",X"22",X"F0",X"22",X"22",X"20",X"00",X"9C",X"99",X"33",X"00",X"2C",X"29",X"00",X"00",
		X"92",X"29",X"22",X"00",X"22",X"22",X"20",X"F0",X"93",X"33",X"02",X"F0",X"C9",X"22",X"20",X"0F",
		X"22",X"29",X"02",X"00",X"CC",X"92",X"20",X"F0",X"92",X"29",X"00",X"00",X"99",X"99",X"FF",X"F0",
		X"00",X"00",X"F0",X"0F",X"00",X"00",X"F2",X"00",X"00",X"00",X"22",X"00",X"00",X"F0",X"22",X"0F",
		X"00",X"00",X"22",X"0F",X"00",X"F0",X"22",X"0F",X"00",X"F0",X"29",X"F0",X"00",X"00",X"92",X"00",
		X"00",X"00",X"22",X"FF",X"00",X"00",X"20",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"CC",X"99",X"99",
		X"00",X"92",X"22",X"99",X"00",X"29",X"22",X"22",X"00",X"92",X"2C",X"22",X"00",X"99",X"99",X"99",
		X"09",X"29",X"29",X"22",X"09",X"99",X"92",X"22",X"09",X"22",X"92",X"22",X"09",X"22",X"99",X"99",
		X"09",X"C2",X"2C",X"99",X"09",X"22",X"C2",X"92",X"09",X"92",X"22",X"22",X"00",X"99",X"29",X"29",
		X"00",X"C2",X"99",X"99",X"00",X"22",X"22",X"92",X"00",X"C2",X"22",X"22",X"00",X"22",X"22",X"C2",
		X"00",X"99",X"99",X"22",X"00",X"CC",X"22",X"9C",X"00",X"CC",X"2C",X"C9",X"00",X"CC",X"22",X"22",
		X"00",X"22",X"22",X"22",X"09",X"99",X"2C",X"29",X"00",X"C9",X"99",X"99",X"00",X"CC",X"22",X"99",
		X"00",X"22",X"2C",X"99",X"00",X"2C",X"22",X"C9",X"00",X"22",X"22",X"C9",X"00",X"22",X"22",X"C9",
		X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"F0",X"99",X"99",X"99",X"00",
		X"22",X"22",X"22",X"90",X"22",X"22",X"22",X"92",X"22",X"22",X"29",X"92",X"99",X"99",X"99",X"29",
		X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"29",X"92",X"99",X"99",X"99",X"00",
		X"99",X"00",X"00",X"02",X"99",X"99",X"00",X"F0",X"22",X"92",X"00",X"F0",X"2C",X"29",X"99",X"00",
		X"22",X"22",X"29",X"FF",X"9C",X"99",X"29",X"00",X"22",X"22",X"92",X"00",X"92",X"29",X"99",X"00",
		X"22",X"92",X"22",X"00",X"99",X"99",X"99",X"00",X"29",X"99",X"2F",X"0F",X"C2",X"22",X"29",X"00",
		X"92",X"C2",X"92",X"0F",X"22",X"9C",X"29",X"00",X"99",X"22",X"20",X"F0",X"99",X"C9",X"92",X"00",
		X"33",X"22",X"29",X"F0",X"33",X"22",X"F9",X"00",X"39",X"92",X"92",X"00",X"33",X"22",X"22",X"F0",
		X"00",X"C9",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"C2",X"22",X"22",
		X"00",X"C2",X"22",X"22",X"00",X"99",X"99",X"99",X"00",X"22",X"99",X"92",X"00",X"22",X"90",X"92",
		X"00",X"22",X"09",X"92",X"00",X"C2",X"90",X"22",X"00",X"C9",X"99",X"99",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"92",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"C2",X"22",X"33",
		X"00",X"C9",X"99",X"29",X"00",X"3C",X"22",X"22",X"00",X"39",X"CC",X"22",X"00",X"39",X"92",X"92",
		X"00",X"39",X"29",X"99",X"00",X"39",X"99",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"20",X"00",
		X"00",X"92",X"00",X"00",X"00",X"29",X"02",X"00",X"00",X"99",X"20",X"00",X"00",X"F0",X"02",X"00",
		X"00",X"00",X"F2",X"00",X"00",X"F0",X"22",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"0F",X"00",
		X"99",X"99",X"09",X"00",X"92",X"29",X"29",X"F0",X"22",X"92",X"92",X"FF",X"29",X"22",X"29",X"F0",
		X"C2",X"92",X"99",X"00",X"C9",X"39",X"02",X"00",X"92",X"92",X"22",X"00",X"22",X"22",X"99",X"00",
		X"92",X"29",X"22",X"00",X"22",X"22",X"99",X"F0",X"9C",X"99",X"29",X"FF",X"2C",X"29",X"90",X"00",
		X"92",X"29",X"22",X"0F",X"22",X"22",X"99",X"0F",X"93",X"33",X"22",X"F0",X"C9",X"22",X"99",X"00",
		X"22",X"29",X"02",X"00",X"CC",X"92",X"20",X"00",X"92",X"29",X"F0",X"0F",X"99",X"99",X"F0",X"F0",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"F0",
		X"00",X"00",X"22",X"0F",X"00",X"00",X"22",X"0F",X"00",X"00",X"29",X"00",X"00",X"00",X"92",X"00",
		X"00",X"00",X"22",X"0F",X"00",X"00",X"20",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"AA",X"00",X"00",X"A6",X"A9",X"00",
		X"00",X"36",X"AA",X"AA",X"00",X"36",X"E9",X"99",X"00",X"A6",X"AA",X"99",X"00",X"3A",X"99",X"99",
		X"00",X"99",X"A9",X"A3",X"00",X"FF",X"A3",X"3A",X"00",X"99",X"97",X"A0",X"00",X"FF",X"AA",X"9F",
		X"00",X"99",X"AA",X"9F",X"00",X"FF",X"9A",X"9F",X"00",X"99",X"59",X"9F",X"00",X"FF",X"E5",X"9F",
		X"00",X"9F",X"AA",X"F5",X"00",X"FF",X"EA",X"FF",X"00",X"99",X"AE",X"FF",X"00",X"AA",X"EA",X"F5",
		X"00",X"69",X"AE",X"F5",X"00",X"F9",X"E5",X"FF",X"00",X"69",X"99",X"FF",X"00",X"EE",X"99",X"3F",
		X"00",X"EE",X"99",X"AF",X"00",X"99",X"A9",X"E3",X"00",X"F5",X"99",X"9E",X"00",X"D9",X"99",X"99",
		X"00",X"00",X"D9",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"99",X"00",
		X"FF",X"99",X"5E",X"00",X"99",X"FF",X"EE",X"90",X"9E",X"99",X"99",X"90",X"EA",X"AA",X"F9",X"90",
		X"EA",X"AA",X"99",X"99",X"AA",X"AA",X"57",X"49",X"EA",X"AA",X"AA",X"A4",X"AA",X"94",X"AA",X"5A",
		X"AA",X"94",X"AA",X"59",X"AA",X"94",X"AA",X"95",X"AA",X"49",X"AA",X"A9",X"EA",X"99",X"AA",X"E9",
		X"AE",X"44",X"AA",X"E9",X"EA",X"99",X"AA",X"59",X"AE",X"99",X"AA",X"59",X"EA",X"44",X"AA",X"59",
		X"EE",X"44",X"A5",X"90",X"EE",X"AE",X"AE",X"90",X"99",X"EA",X"E5",X"90",X"F9",X"EE",X"E5",X"90",
		X"99",X"99",X"59",X"50",X"99",X"F9",X"99",X"90",X"D9",X"99",X"99",X"90",X"00",X"9A",X"99",X"40",
		X"00",X"99",X"39",X"0F",X"00",X"09",X"99",X"0F",X"00",X"00",X"99",X"F0",X"00",X"00",X"00",X"F0",
		X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"AE",X"E9",X"00",
		X"00",X"9A",X"AE",X"00",X"00",X"F9",X"99",X"99",X"00",X"FF",X"A9",X"AE",X"00",X"99",X"99",X"9A",
		X"00",X"9A",X"99",X"A9",X"00",X"9A",X"97",X"A9",X"00",X"9A",X"95",X"99",X"00",X"99",X"A5",X"A7",
		X"00",X"99",X"A5",X"EA",X"05",X"EE",X"E5",X"AE",X"05",X"EE",X"E5",X"EA",X"05",X"EE",X"E5",X"AE",
		X"05",X"EE",X"5E",X"EA",X"05",X"9E",X"55",X"EE",X"05",X"9E",X"5E",X"EE",X"53",X"9E",X"55",X"EE",
		X"55",X"A9",X"65",X"EE",X"05",X"5A",X"AA",X"E5",X"05",X"EE",X"DD",X"65",X"05",X"55",X"DD",X"AA",
		X"05",X"EE",X"DD",X"DD",X"00",X"0E",X"AA",X"FF",X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"9A",X"95",X"00",X"00",X"A9",X"95",X"00",X"00",
		X"99",X"59",X"00",X"00",X"A7",X"59",X"00",X"00",X"AA",X"59",X"00",X"00",X"A7",X"59",X"00",X"00",
		X"AA",X"59",X"00",X"00",X"A7",X"59",X"00",X"00",X"AA",X"59",X"00",X"00",X"A7",X"59",X"00",X"00",
		X"A9",X"59",X"00",X"00",X"79",X"59",X"00",X"00",X"A9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"DA",X"99",X"00",X"00",X"DD",X"90",X"00",X"00",
		X"DD",X"99",X"00",X"00",X"AA",X"90",X"00",X"00",X"AE",X"90",X"00",X"00",X"E9",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"EA",X"00",X"EE",
		X"05",X"EE",X"99",X"EE",X"05",X"5A",X"EA",X"99",X"05",X"EE",X"A9",X"A9",X"55",X"AA",X"9A",X"FF",
		X"53",X"99",X"A9",X"A9",X"59",X"7A",X"99",X"99",X"59",X"AA",X"A7",X"A7",X"5F",X"AA",X"EA",X"EA",
		X"59",X"AA",X"5E",X"AE",X"59",X"A9",X"EE",X"EA",X"5F",X"99",X"5E",X"AE",X"59",X"99",X"EE",X"EA",
		X"59",X"39",X"5E",X"EE",X"5F",X"E9",X"E5",X"EA",X"59",X"E9",X"5E",X"EE",X"59",X"EE",X"E5",X"EE",
		X"5F",X"EE",X"5E",X"5E",X"59",X"EE",X"56",X"65",X"59",X"E5",X"AA",X"AA",X"53",X"99",X"DD",X"DD",
		X"55",X"AA",X"DD",X"FF",X"05",X"5E",X"DD",X"DD",X"05",X"E5",X"AA",X"AA",X"05",X"5E",X"EE",X"AE",
		X"05",X"EE",X"90",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",
		X"AE",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"A9",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"97",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"DA",X"99",X"00",X"00",
		X"DD",X"90",X"00",X"00",X"DD",X"90",X"00",X"00",X"AA",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",
		X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"A9",X"00",
		X"00",X"5E",X"AA",X"99",X"00",X"E9",X"99",X"AA",X"00",X"99",X"99",X"EE",X"09",X"99",X"3F",X"55",
		X"09",X"94",X"35",X"55",X"09",X"43",X"55",X"99",X"09",X"49",X"FF",X"BA",X"95",X"94",X"FF",X"EE",
		X"99",X"AA",X"FF",X"EE",X"95",X"A4",X"FF",X"EE",X"99",X"49",X"FF",X"EE",X"95",X"94",X"FF",X"EE",
		X"99",X"74",X"FF",X"EE",X"09",X"EE",X"55",X"EE",X"09",X"99",X"55",X"EE",X"00",X"99",X"55",X"EE",
		X"00",X"EA",X"5F",X"3B",X"00",X"AA",X"F5",X"99",X"00",X"EE",X"33",X"53",X"00",X"9E",X"9E",X"53",
		X"00",X"09",X"AE",X"E3",X"00",X"00",X"99",X"A3",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"3A",X"99",X"00",X"00",X"33",X"34",X"00",X"00",
		X"99",X"40",X"00",X"00",X"55",X"40",X"00",X"00",X"9C",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"B5",X"30",X"00",X"00",X"55",X"00",X"00",X"00",
		X"FF",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"55",X"90",X"00",X"00",
		X"55",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"5E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9A",X"00",X"00",X"99",X"A3",X"00",X"09",X"AE",X"E3",
		X"00",X"9E",X"9E",X"53",X"00",X"EE",X"33",X"53",X"00",X"EE",X"F5",X"99",X"00",X"EA",X"5F",X"3B",
		X"00",X"99",X"55",X"EE",X"09",X"99",X"55",X"EE",X"09",X"EE",X"55",X"EE",X"99",X"74",X"FF",X"EE",
		X"95",X"94",X"FF",X"EE",X"99",X"49",X"FF",X"EE",X"95",X"A4",X"FF",X"EE",X"99",X"AA",X"FF",X"EE",
		X"95",X"94",X"FF",X"EE",X"09",X"49",X"FF",X"BA",X"09",X"43",X"55",X"99",X"09",X"94",X"35",X"55",
		X"09",X"99",X"3F",X"55",X"00",X"99",X"99",X"EE",X"00",X"E9",X"99",X"AA",X"00",X"AA",X"AA",X"99",
		X"00",X"EE",X"A9",X"00",X"00",X"EE",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"55",X"90",X"00",X"00",
		X"55",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"55",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",
		X"55",X"00",X"00",X"00",X"B5",X"30",X"00",X"00",X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"9C",X"00",X"00",X"00",X"55",X"40",X"00",X"00",X"99",X"40",X"00",X"00",
		X"93",X"94",X"00",X"00",X"3A",X"99",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"90",X"90",X"99",X"00",X"09",X"09",X"99",X"00",X"99",X"90",X"22",
		X"00",X"99",X"99",X"22",X"92",X"33",X"99",X"22",X"FF",X"A3",X"99",X"22",X"F3",X"3A",X"22",X"22",
		X"F2",X"A3",X"92",X"22",X"09",X"99",X"29",X"22",X"93",X"33",X"29",X"22",X"92",X"95",X"29",X"22",
		X"99",X"55",X"29",X"22",X"9F",X"55",X"29",X"22",X"99",X"55",X"29",X"22",X"9F",X"55",X"29",X"22",
		X"99",X"99",X"69",X"22",X"9F",X"FF",X"29",X"22",X"99",X"FF",X"29",X"22",X"9F",X"FF",X"29",X"22",
		X"99",X"1F",X"29",X"22",X"92",X"1F",X"29",X"22",X"93",X"33",X"29",X"22",X"09",X"93",X"29",X"22",
		X"F2",X"A3",X"02",X"22",X"F2",X"3A",X"22",X"22",X"F2",X"A3",X"00",X"22",X"92",X"33",X"00",X"22",
		X"00",X"90",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"22",X"00",X"00",X"55",X"11",X"00",X"00",X"55",X"11",X"00",X"00",X"55",X"15",
		X"00",X"55",X"55",X"15",X"00",X"55",X"55",X"15",X"00",X"55",X"55",X"53",X"00",X"55",X"11",X"33",
		X"00",X"53",X"11",X"17",X"00",X"14",X"33",X"99",X"99",X"41",X"33",X"BB",X"00",X"11",X"3A",X"99",
		X"00",X"55",X"A9",X"99",X"00",X"55",X"AB",X"29",X"00",X"55",X"AB",X"32",X"00",X"55",X"AB",X"22",
		X"00",X"FF",X"AB",X"22",X"00",X"FF",X"AB",X"55",X"00",X"FF",X"AB",X"59",X"00",X"FF",X"A9",X"99",
		X"00",X"11",X"5A",X"99",X"99",X"41",X"FF",X"BB",X"00",X"11",X"FF",X"FF",X"00",X"55",X"11",X"11",
		X"00",X"55",X"51",X"55",X"00",X"55",X"55",X"55",X"00",X"FF",X"55",X"35",X"00",X"FF",X"55",X"1F",
		X"00",X"00",X"FF",X"19",X"00",X"00",X"FF",X"11",X"00",X"00",X"FF",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"90",X"F0",X"00",X"00",X"59",X"00",X"00",X"00",
		X"55",X"39",X"00",X"00",X"95",X"99",X"00",X"00",X"11",X"F9",X"00",X"00",X"11",X"11",X"30",X"00",
		X"99",X"99",X"F0",X"00",X"99",X"FF",X"00",X"00",X"59",X"99",X"00",X"00",X"59",X"FF",X"00",X"00",
		X"59",X"FF",X"00",X"00",X"59",X"99",X"00",X"00",X"99",X"FF",X"00",X"00",X"99",X"99",X"F0",X"00",
		X"44",X"11",X"00",X"00",X"11",X"FF",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"F9",X"00",X"00",
		X"50",X"0F",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EE",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"EE",X"00",X"00",X"99",X"99",X"00",X"00",
		X"22",X"92",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"09",X"00",
		X"99",X"99",X"00",X"00",X"92",X"33",X"09",X"00",X"22",X"33",X"00",X"00",X"22",X"99",X"F9",X"00",
		X"22",X"99",X"F0",X"09",X"22",X"33",X"F9",X"99",X"22",X"33",X"F9",X"99",X"29",X"99",X"3F",X"99",
		X"22",X"29",X"3F",X"99",X"22",X"22",X"FF",X"90",X"22",X"22",X"F3",X"90",X"22",X"22",X"F3",X"00",
		X"29",X"99",X"F9",X"00",X"22",X"22",X"F9",X"00",X"22",X"22",X"F9",X"00",X"22",X"22",X"99",X"00",
		X"22",X"22",X"99",X"00",X"22",X"22",X"99",X"00",X"29",X"92",X"99",X"00",X"22",X"22",X"99",X"00",
		X"22",X"22",X"99",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"9F",X"00",X"22",X"22",X"FF",X"00",
		X"11",X"11",X"FF",X"00",X"11",X"11",X"9F",X"00",X"11",X"11",X"99",X"00",X"11",X"11",X"99",X"00",
		X"11",X"11",X"99",X"00",X"11",X"11",X"99",X"00",X"22",X"22",X"99",X"00",X"21",X"22",X"99",X"00",
		X"21",X"22",X"99",X"00",X"21",X"91",X"F9",X"00",X"21",X"11",X"F9",X"00",X"91",X"11",X"F9",X"00",
		X"92",X"11",X"F3",X"00",X"92",X"11",X"F3",X"90",X"92",X"22",X"FF",X"90",X"92",X"19",X"3F",X"99",
		X"99",X"99",X"3F",X"99",X"92",X"33",X"F9",X"99",X"92",X"33",X"F9",X"99",X"92",X"99",X"F0",X"09",
		X"92",X"99",X"F9",X"00",X"11",X"33",X"00",X"00",X"22",X"33",X"09",X"00",X"11",X"99",X"00",X"00",
		X"11",X"99",X"09",X"00",X"11",X"99",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"91",X"00",X"00",
		X"99",X"99",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"99",X"00",X"00",X"EE",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"15",X"00",X"00",
		X"90",X"15",X"50",X"00",X"99",X"F1",X"55",X"00",X"99",X"11",X"55",X"00",X"F9",X"11",X"55",X"00",
		X"F9",X"11",X"55",X"00",X"F5",X"55",X"55",X"00",X"FF",X"55",X"55",X"00",X"FF",X"55",X"55",X"00",
		X"FF",X"F5",X"15",X"50",X"FF",X"FF",X"11",X"55",X"0F",X"F3",X"11",X"55",X"0F",X"F3",X"11",X"55",
		X"0F",X"F3",X"31",X"11",X"0F",X"F3",X"5F",X"11",X"0F",X"F3",X"9F",X"19",X"00",X"FF",X"BB",X"99",
		X"00",X"1F",X"9B",X"99",X"00",X"1F",X"99",X"59",X"00",X"11",X"99",X"55",X"00",X"11",X"91",X"25",
		X"00",X"11",X"51",X"25",X"00",X"11",X"51",X"25",X"00",X"51",X"55",X"22",X"00",X"51",X"95",X"22",
		X"00",X"51",X"99",X"12",X"00",X"51",X"B9",X"91",X"00",X"51",X"BB",X"33",X"00",X"51",X"FB",X"F3",
		X"55",X"11",X"5F",X"99",X"05",X"51",X"FF",X"99",X"05",X"55",X"FF",X"FF",X"00",X"F5",X"3F",X"F0",
		X"00",X"0F",X"9F",X"FF",X"00",X"00",X"99",X"19",X"00",X"99",X"19",X"99",X"00",X"09",X"11",X"3F",
		X"00",X"00",X"F1",X"31",X"00",X"00",X"F1",X"99",X"00",X"00",X"9F",X"F9",X"00",X"00",X"90",X"FF",
		X"00",X"00",X"90",X"FF",X"00",X"00",X"90",X"FF",X"00",X"00",X"90",X"FF",X"00",X"00",X"90",X"FF",
		X"00",X"00",X"99",X"3F",X"00",X"00",X"99",X"39",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"09",
		X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"33",X"90",X"90",X"00",X"55",X"99",X"00",X"00",X"15",X"33",X"00",
		X"00",X"11",X"FF",X"90",X"01",X"11",X"5F",X"99",X"01",X"11",X"55",X"33",X"90",X"55",X"55",X"5F",
		X"99",X"55",X"15",X"FF",X"19",X"55",X"11",X"5F",X"F1",X"55",X"11",X"11",X"51",X"55",X"51",X"11",
		X"05",X"FF",X"F9",X"11",X"0F",X"FF",X"5F",X"11",X"00",X"FF",X"F9",X"11",X"00",X"1F",X"99",X"11",
		X"00",X"11",X"99",X"F1",X"00",X"11",X"9B",X"BB",X"00",X"51",X"9B",X"99",X"00",X"55",X"9B",X"29",
		X"00",X"55",X"BB",X"22",X"00",X"55",X"FB",X"12",X"00",X"55",X"11",X"19",X"00",X"FF",X"11",X"99",
		X"00",X"FF",X"11",X"9D",X"00",X"FF",X"11",X"FD",X"00",X"FF",X"21",X"1D",X"00",X"0F",X"51",X"11",
		X"00",X"00",X"51",X"55",X"00",X"00",X"51",X"F5",X"00",X"00",X"52",X"FF",X"00",X"00",X"FF",X"FF",
		X"11",X"FF",X"99",X"00",X"11",X"55",X"99",X"00",X"11",X"55",X"11",X"00",X"FF",X"55",X"19",X"00",
		X"99",X"11",X"99",X"00",X"99",X"11",X"99",X"00",X"9F",X"11",X"99",X"00",X"5F",X"F1",X"33",X"00",
		X"5F",X"BB",X"53",X"00",X"95",X"99",X"5F",X"09",X"9F",X"99",X"55",X"00",X"FF",X"99",X"55",X"09",
		X"FF",X"92",X"15",X"00",X"11",X"95",X"15",X"99",X"11",X"95",X"19",X"FF",X"11",X"99",X"F1",X"00",
		X"51",X"B9",X"99",X"00",X"55",X"1F",X"99",X"99",X"55",X"11",X"99",X"F9",X"5F",X"91",X"9F",X"9F",
		X"55",X"95",X"9F",X"19",X"FF",X"95",X"19",X"91",X"FF",X"95",X"11",X"55",X"FF",X"95",X"55",X"55",
		X"FF",X"99",X"55",X"55",X"00",X"99",X"00",X"95",X"00",X"90",X"00",X"19",X"00",X"00",X"00",X"11",
		X"00",X"00",X"90",X"F1",X"00",X"00",X"F9",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"C9",X"99",X"90",X"00",X"BC",X"99",X"99",
		X"00",X"B6",X"99",X"99",X"00",X"AA",X"9C",X"99",X"00",X"AC",X"C0",X"99",X"00",X"AA",X"BE",X"99",
		X"04",X"EA",X"BB",X"CB",X"04",X"BB",X"BA",X"E9",X"00",X"EE",X"BE",X"0C",X"00",X"BB",X"5B",X"CB",
		X"00",X"EB",X"BB",X"E0",X"00",X"FE",X"5B",X"BC",X"00",X"B5",X"BB",X"BB",X"04",X"BB",X"F5",X"BE",
		X"4C",X"BB",X"B5",X"BB",X"50",X"BB",X"5B",X"BB",X"50",X"BB",X"B5",X"BB",X"00",X"66",X"5B",X"BB",
		X"00",X"BB",X"BF",X"BB",X"00",X"9C",X"FB",X"BB",X"00",X"EB",X"BB",X"69",X"00",X"BE",X"6F",X"9B",
		X"00",X"C9",X"BB",X"BB",X"00",X"00",X"00",X"BC",X"00",X"00",X"CC",X"C9",X"00",X"00",X"00",X"9B",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"99",
		X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"9A",X"00",X"99",X"CC",X"C9",X"00",X"99",X"00",X"BC",
		X"00",X"C9",X"AB",X"AB",X"00",X"BE",X"BB",X"BB",X"00",X"EB",X"AA",X"B9",X"00",X"9C",X"BB",X"BB",
		X"00",X"AA",X"BB",X"BB",X"00",X"AA",X"BB",X"BB",X"50",X"BB",X"BB",X"BB",X"50",X"BB",X"BB",X"BB",
		X"4C",X"BB",X"B5",X"BB",X"04",X"BB",X"5B",X"BE",X"00",X"BE",X"B5",X"BB",X"00",X"E5",X"5B",X"5C",
		X"00",X"FB",X"55",X"55",X"00",X"BB",X"5B",X"55",X"00",X"EE",X"55",X"0C",X"04",X"BB",X"5A",X"E9",
		X"04",X"EF",X"BB",X"CB",X"00",X"6B",X"BE",X"AA",X"00",X"BB",X"C0",X"00",X"00",X"AA",X"9C",X"00",
		X"00",X"B6",X"AA",X"00",X"00",X"BC",X"00",X"00",X"00",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"D9",X"00",X"00",X"D9",X"99",
		X"00",X"D9",X"99",X"99",X"00",X"F5",X"99",X"9E",X"00",X"99",X"A9",X"E3",X"00",X"EE",X"99",X"AF",
		X"00",X"EE",X"99",X"3F",X"00",X"69",X"99",X"FF",X"00",X"F9",X"E5",X"FF",X"00",X"69",X"AE",X"F5",
		X"00",X"AA",X"EA",X"F5",X"00",X"99",X"AE",X"FF",X"00",X"FF",X"EA",X"FF",X"00",X"9F",X"AA",X"F5",
		X"00",X"FF",X"E5",X"9F",X"00",X"99",X"59",X"9F",X"00",X"FF",X"9A",X"9F",X"00",X"99",X"AA",X"9F",
		X"00",X"FF",X"AA",X"9F",X"00",X"99",X"97",X"A0",X"00",X"FF",X"A3",X"3A",X"00",X"99",X"A9",X"A3",
		X"00",X"3A",X"99",X"99",X"00",X"A6",X"AA",X"99",X"00",X"36",X"E9",X"99",X"00",X"36",X"AA",X"AA",
		X"00",X"A6",X"A9",X"00",X"00",X"9A",X"AA",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"99",X"F0",X"00",X"09",X"99",X"0F",X"00",X"99",X"39",X"0F",
		X"00",X"9A",X"99",X"40",X"D9",X"99",X"99",X"90",X"99",X"F9",X"99",X"90",X"99",X"99",X"59",X"50",
		X"F9",X"EE",X"E5",X"90",X"99",X"EA",X"E5",X"90",X"EE",X"AE",X"AE",X"90",X"EE",X"44",X"A5",X"90",
		X"EA",X"44",X"AA",X"59",X"AE",X"99",X"AA",X"59",X"EA",X"99",X"AA",X"59",X"AE",X"44",X"AA",X"E9",
		X"EA",X"99",X"AA",X"E9",X"AA",X"49",X"AA",X"A9",X"AA",X"94",X"AA",X"95",X"AA",X"94",X"AA",X"59",
		X"AA",X"94",X"AA",X"5A",X"EA",X"AA",X"AA",X"A4",X"AA",X"AA",X"57",X"49",X"EA",X"AA",X"99",X"99",
		X"EA",X"AA",X"F9",X"90",X"9E",X"99",X"99",X"90",X"99",X"FF",X"EE",X"90",X"FF",X"99",X"5E",X"00",
		X"99",X"99",X"99",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"99",X"90",
		X"00",X"DD",X"29",X"99",X"00",X"11",X"22",X"22",X"00",X"11",X"92",X"22",X"00",X"F7",X"19",X"22",
		X"09",X"11",X"93",X"11",X"09",X"11",X"11",X"11",X"09",X"DD",X"1D",X"11",X"09",X"44",X"1D",X"77",
		X"09",X"44",X"17",X"77",X"09",X"44",X"1D",X"77",X"09",X"44",X"17",X"77",X"09",X"45",X"17",X"77",
		X"9F",X"71",X"75",X"77",X"92",X"11",X"F7",X"77",X"92",X"71",X"75",X"77",X"96",X"11",X"F7",X"77",
		X"9F",X"11",X"FF",X"77",X"99",X"77",X"11",X"F7",X"09",X"F2",X"33",X"1F",X"00",X"22",X"99",X"11",
		X"00",X"92",X"22",X"33",X"00",X"09",X"52",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"25",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"09",X"00",X"00",
		X"2A",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",
		X"00",X"00",X"90",X"22",X"00",X"90",X"99",X"22",X"00",X"99",X"22",X"99",X"00",X"92",X"22",X"33",
		X"00",X"22",X"99",X"11",X"09",X"42",X"33",X"17",X"99",X"77",X"11",X"77",X"9F",X"11",X"D7",X"77",
		X"96",X"11",X"DD",X"77",X"92",X"71",X"D7",X"77",X"92",X"14",X"57",X"77",X"9F",X"44",X"77",X"77",
		X"09",X"44",X"15",X"77",X"09",X"44",X"17",X"77",X"09",X"44",X"15",X"77",X"09",X"44",X"15",X"75",
		X"09",X"44",X"1D",X"77",X"09",X"77",X"15",X"11",X"09",X"11",X"11",X"11",X"09",X"11",X"93",X"11",
		X"00",X"F7",X"19",X"22",X"00",X"11",X"92",X"52",X"00",X"11",X"22",X"22",X"00",X"DD",X"59",X"00",
		X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"F9",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",
		X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"25",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"59",X"90",X"00",X"00",X"55",X"99",X"00",X"00",X"05",X"95",X"00",X"00",X"00",X"95",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"95",X"00",
		X"00",X"05",X"95",X"00",X"00",X"55",X"90",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"9A",X"9A",X"00",X"0B",X"AB",X"9B",X"00",X"05",X"BD",X"9D",X"00",X"0F",X"BB",X"9B",
		X"00",X"05",X"5B",X"5B",X"00",X"95",X"BA",X"9A",X"00",X"DD",X"99",X"EE",X"00",X"99",X"EE",X"99",
		X"00",X"DD",X"9E",X"55",X"00",X"99",X"9E",X"99",X"00",X"DD",X"9E",X"9E",X"00",X"99",X"EE",X"59",
		X"00",X"DD",X"E5",X"55",X"0A",X"99",X"EB",X"55",X"0D",X"DD",X"E5",X"55",X"09",X"99",X"EB",X"55",
		X"0A",X"AA",X"B5",X"55",X"0A",X"AB",X"BB",X"55",X"00",X"BA",X"B5",X"55",X"00",X"AB",X"BB",X"55",
		X"00",X"BA",X"BB",X"59",X"00",X"AB",X"A5",X"9F",X"00",X"BA",X"9B",X"99",X"00",X"AB",X"9B",X"F5",
		X"00",X"BA",X"B5",X"59",X"00",X"AB",X"55",X"55",X"00",X"B9",X"99",X"99",X"00",X"0A",X"BA",X"9A",
		X"00",X"0B",X"AB",X"AB",X"00",X"05",X"BB",X"9B",X"00",X"0F",X"B5",X"95",X"00",X"05",X"AB",X"AB",
		X"09",X"99",X"99",X"00",X"9B",X"AB",X"AB",X"00",X"95",X"BD",X"BD",X"00",X"95",X"BB",X"BB",X"00",
		X"95",X"5B",X"5B",X"00",X"95",X"BA",X"BA",X"00",X"EE",X"DD",X"55",X"00",X"99",X"DD",X"DD",X"00",
		X"59",X"BB",X"BB",X"00",X"9E",X"DD",X"DD",X"00",X"59",X"BB",X"BB",X"00",X"EA",X"DD",X"DD",X"00",
		X"59",X"BB",X"BB",X"00",X"EA",X"DB",X"DB",X"00",X"E9",X"BB",X"BB",X"00",X"59",X"BB",X"BB",X"00",
		X"EA",X"BA",X"BB",X"00",X"59",X"BB",X"BB",X"00",X"E9",X"AB",X"AB",X"00",X"E9",X"BB",X"BB",X"00",
		X"59",X"AA",X"AA",X"00",X"59",X"BB",X"BB",X"00",X"59",X"AA",X"AA",X"00",X"55",X"B9",X"99",X"00",
		X"55",X"AA",X"C5",X"00",X"55",X"B9",X"9B",X"00",X"99",X"99",X"99",X"00",X"BB",X"AB",X"AB",X"00",
		X"A5",X"BA",X"BA",X"00",X"A5",X"BB",X"BB",X"00",X"05",X"B5",X"BB",X"00",X"05",X"AB",X"AB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"FB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"00",X"BF",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"FB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"B0",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"FB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"BB",X"FF",X"BB",
		X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BF",X"0B",X"BB",X"00",X"FB",X"00",X"BF",
		X"00",X"BB",X"00",X"BB",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"FB",X"00",X"00",X"BB",X"FB",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"FF",X"00",X"BB",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"FF",X"0B",X"00",X"00",X"FF",X"BB",X"BB",
		X"00",X"FF",X"BB",X"FB",X"00",X"BF",X"BB",X"FF",X"00",X"BF",X"BB",X"BF",X"00",X"BF",X"BB",X"BB",
		X"00",X"BF",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"B0",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"BF",X"BB",X"FF",
		X"00",X"BB",X"BB",X"FF",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"00",X"BB",
		X"00",X"BB",X"00",X"BB",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FB",X"00",X"00",X"BB",X"FB",X"00",
		X"00",X"BB",X"FB",X"00",X"00",X"BB",X"FB",X"00",X"00",X"BB",X"FB",X"00",X"00",X"BB",X"FB",X"00",
		X"00",X"FF",X"BB",X"00",X"00",X"BF",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BF",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"BB",
		X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BF",X"BB",X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"FF",X"BB",X"00",X"FB",X"FB",X"BB",
		X"00",X"FB",X"BB",X"BB",X"00",X"FB",X"BB",X"BB",X"00",X"FB",X"BB",X"BB",X"00",X"FF",X"BB",X"FB",
		X"00",X"FF",X"BB",X"FB",X"00",X"FF",X"BB",X"FF",X"00",X"FF",X"BB",X"FF",X"00",X"BF",X"BB",X"FF",
		X"00",X"BB",X"BB",X"FF",X"00",X"BB",X"BB",X"FF",X"00",X"BB",X"BB",X"FF",X"00",X"BB",X"B0",X"BF",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"BB",X"BF",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"FF",X"BB",X"FF",X"00",X"FB",X"0B",X"BB",X"00",X"BB",X"00",X"BB",
		X"00",X"BB",X"00",X"BB",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"FF",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FB",X"00",
		X"00",X"BB",X"FB",X"00",X"00",X"BB",X"FB",X"00",X"00",X"BB",X"FB",X"00",X"00",X"FB",X"BB",X"00",
		X"00",X"FB",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"FF",X"BB",X"B0",X"00",X"FF",X"BB",X"BB",
		X"00",X"FF",X"BB",X"BB",X"00",X"BB",X"FF",X"BB",X"00",X"00",X"BF",X"BB",X"00",X"00",X"BB",X"FB",
		X"00",X"B0",X"00",X"BF",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"FB",X"00",X"BB",X"BB",X"FB",X"00",X"BB",X"BB",X"FB",
		X"00",X"FB",X"BB",X"FB",X"00",X"FF",X"BB",X"FF",X"00",X"FF",X"BB",X"FF",X"00",X"FF",X"B0",X"FF",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"BB",X"FB",X"BB",
		X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BF",X"0B",X"FB",X"00",X"FF",X"00",X"FF",
		X"00",X"FB",X"00",X"BB",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"11",X"11",X"10",X"00",X"11",X"11",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"01",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"10",
		X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"01",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"01",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"10",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"11",X"00",X"11",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",
		X"00",X"11",X"11",X"10",X"00",X"11",X"11",X"10",X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"10",
		X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"10",X"00",X"11",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"EE",X"A0",X"00",X"00",X"23",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"00",X"5E",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"E0",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"33",X"A0",X"00",X"00",X"53",X"A0",
		X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"53",X"00",
		X"00",X"00",X"23",X"A0",X"00",X"00",X"33",X"00",X"00",X"00",X"0E",X"A0",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"E0",X"A0",X"00",X"00",X"EE",X"A0",X"00",X"00",X"33",X"00",X"00",X"00",X"23",X"00",
		X"00",X"00",X"23",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"EE",X"A0",X"00",X"00",X"E0",X"A0",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"F9",X"F0",X"00",X"00",X"99",X"F5",X"00",X"00",X"99",X"9B",
		X"00",X"00",X"99",X"9F",X"00",X"00",X"09",X"95",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"09",X"09",X"00",X"99",X"99",X"99",
		X"00",X"FF",X"99",X"05",X"00",X"EE",X"EE",X"EE",X"00",X"BB",X"BB",X"BB",X"0E",X"44",X"99",X"F5",
		X"0F",X"77",X"59",X"F9",X"5F",X"55",X"55",X"99",X"59",X"55",X"9F",X"55",X"59",X"FF",X"5F",X"FF",
		X"59",X"B5",X"FF",X"FF",X"5F",X"5E",X"FF",X"FF",X"5F",X"55",X"FF",X"FF",X"5F",X"55",X"FF",X"FF",
		X"5F",X"F5",X"FF",X"FF",X"5F",X"FF",X"FF",X"FF",X"5F",X"FF",X"FF",X"FF",X"59",X"FF",X"FF",X"FF",
		X"59",X"55",X"5F",X"FF",X"59",X"55",X"9F",X"55",X"5F",X"55",X"55",X"99",X"0F",X"77",X"F9",X"F9",
		X"0E",X"44",X"99",X"F5",X"00",X"BB",X"BB",X"BB",X"00",X"FF",X"FF",X"EF",X"00",X"FF",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"E9",X"90",X"00",X"00",X"B9",X"99",X"00",X"00",X"9F",X"90",X"00",X"00",
		X"0F",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",X"FE",X"99",X"00",X"00",
		X"FE",X"59",X"00",X"00",X"FE",X"59",X"00",X"00",X"FE",X"59",X"00",X"00",X"FE",X"99",X"00",X"00",
		X"FE",X"99",X"00",X"00",X"FE",X"59",X"00",X"00",X"FE",X"59",X"00",X"00",X"FE",X"59",X"00",X"00",
		X"FE",X"90",X"00",X"00",X"FF",X"09",X"00",X"00",X"5F",X"90",X"00",X"00",X"95",X"00",X"00",X"00",
		X"9F",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
