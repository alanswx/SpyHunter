library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_cpu is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(15 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_cpu is
	type rom is array(0 to  57343) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"00",X"01",X"5D",X"C4",X"4B",X"4C",X"19",X"2B",X"02",X"3D",X"02",X"10",X"00",X"AF",X"01",
		X"18",X"FE",X"39",X"C0",X"CA",X"41",X"CF",X"D0",X"53",X"99",X"5B",X"03",X"8F",X"97",X"9C",X"1A",
		X"DF",X"5C",X"39",X"D4",X"4A",X"3C",X"07",X"4C",X"18",X"82",X"28",X"C4",X"17",X"E1",X"17",X"C5",
		X"48",X"85",X"D1",X"4F",X"52",X"0B",X"D7",X"81",X"80",X"5A",X"A8",X"05",X"D9",X"54",X"9C",X"08",
		X"E5",X"B8",X"7A",X"D3",X"E9",X"89",X"DE",X"1A",X"72",X"0C",X"7B",X"DB",X"89",X"F5",X"9A",X"3B",
		X"89",X"EF",X"29",X"4F",X"7B",X"0F",X"C2",X"81",X"EB",X"4A",X"EB",X"42",X"8B",X"A9",X"D2",X"73",
		X"2E",X"FB",X"29",X"B8",X"6E",X"E3",X"3E",X"07",X"D3",X"E8",X"76",X"43",X"4F",X"50",X"59",X"52",
		X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"32",X"20",X"42",X"41",X"4C",X"4C",X"59",X"20",
		X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"4D",X"46",X"47",X"20",X"43",X"4F",X"00",X"00",X"00",
		X"00",X"12",X"8C",X"52",X"82",X"64",X"74",X"B7",X"16",X"91",X"9D",X"83",X"AB",X"86",X"A1",X"C2",
		X"72",X"BB",X"84",X"91",X"FA",X"93",X"95",X"F7",X"10",X"94",X"C7",X"B4",X"08",X"FA",X"64",X"4D",
		X"CD",X"02",X"36",X"F6",X"19",X"0B",X"7D",X"C4",X"FA",X"56",X"F1",X"E4",X"8F",X"4E",X"4D",X"87",
		X"A8",X"ED",X"AE",X"B3",X"EE",X"FB",X"71",X"39",X"BD",X"20",X"DA",X"F2",X"B4",X"E4",X"31",X"F1",
		X"E7",X"E5",X"FA",X"EA",X"B5",X"B7",X"EA",X"70",X"9D",X"0C",X"B3",X"A8",X"E4",X"A9",X"7A",X"0B",
		X"97",X"7A",X"29",X"33",X"CB",X"FB",X"E0",X"65",X"8E",X"2F",X"22",X"B1",X"AF",X"EC",X"38",X"78",
		X"EE",X"E6",X"A9",X"0D",X"62",X"CE",X"D8",X"32",X"66",X"E7",X"4F",X"A7",X"FE",X"28",X"E2",X"73",
		X"F3",X"21",X"64",X"00",X"2B",X"7C",X"B5",X"20",X"FB",X"D3",X"E0",X"AF",X"D3",X"00",X"3E",X"02",
		X"D3",X"E8",X"06",X"09",X"AF",X"D3",X"E8",X"3C",X"D3",X"E8",X"10",X"F8",X"3E",X"05",X"D3",X"E8",
		X"31",X"FE",X"F7",X"CD",X"5D",X"0A",X"CD",X"B6",X"07",X"28",X"04",X"D3",X"E0",X"18",X"FC",X"CD",
		X"2B",X"3D",X"3E",X"01",X"32",X"16",X"F4",X"CD",X"26",X"13",X"3E",X"55",X"32",X"00",X"F4",X"ED",
		X"5E",X"3E",X"00",X"ED",X"47",X"3E",X"08",X"D3",X"F0",X"3E",X"C7",X"D3",X"F3",X"3E",X"01",X"D3",
		X"F3",X"3E",X"A7",X"D3",X"F1",X"3E",X"9C",X"D3",X"F1",X"3E",X"01",X"32",X"13",X"F4",X"3E",X"02",
		X"32",X"14",X"F4",X"3E",X"40",X"32",X"15",X"F4",X"CD",X"93",X"01",X"21",X"1E",X"F4",X"22",X"1B",
		X"F4",X"FB",X"CD",X"85",X"0B",X"CD",X"F9",X"3C",X"0E",X"02",X"CD",X"4E",X"3D",X"CD",X"F9",X"3C",
		X"CD",X"F9",X"3C",X"0E",X"02",X"CD",X"4E",X"3D",X"0E",X"01",X"CD",X"4E",X"3D",X"CD",X"F9",X"3C",
		X"C3",X"0F",X"89",X"06",X"20",X"21",X"FF",X"EB",X"36",X"5B",X"2B",X"10",X"FB",X"01",X"C0",X"03",
		X"36",X"00",X"E5",X"D1",X"1B",X"ED",X"B8",X"06",X"20",X"36",X"5B",X"2B",X"10",X"FB",X"C9",X"08",
		X"D9",X"DD",X"E5",X"FD",X"E5",X"AF",X"32",X"04",X"F4",X"3E",X"A7",X"D3",X"F0",X"3E",X"18",X"D3",
		X"F0",X"CD",X"16",X"05",X"CD",X"31",X"06",X"CD",X"E3",X"06",X"3A",X"8A",X"F3",X"B7",X"28",X"1D",
		X"21",X"8D",X"F3",X"7E",X"D6",X"01",X"77",X"F2",X"EC",X"01",X"36",X"1E",X"2B",X"7E",X"C6",X"01",
		X"27",X"FE",X"60",X"20",X"07",X"36",X"00",X"2B",X"7E",X"C6",X"01",X"27",X"77",X"2A",X"91",X"F0",
		X"7D",X"D3",X"84",X"7C",X"D3",X"85",X"3A",X"0A",X"F0",X"B7",X"28",X"1F",X"CB",X"7F",X"3E",X"FF",
		X"28",X"01",X"AF",X"21",X"0D",X"F0",X"BE",X"20",X"0F",X"B7",X"28",X"05",X"3E",X"20",X"32",X"38",
		X"F0",X"AF",X"32",X"0A",X"F0",X"32",X"0C",X"F0",X"7E",X"D3",X"86",X"FB",X"3A",X"04",X"F4",X"B7",
		X"28",X"FA",X"FD",X"E1",X"DD",X"E1",X"D9",X"08",X"FB",X"ED",X"4D",X"F5",X"3A",X"8F",X"F3",X"3C",
		X"32",X"8F",X"F3",X"3E",X"03",X"D3",X"F0",X"32",X"04",X"F4",X"F1",X"ED",X"4D",X"F5",X"E5",X"C5",
		X"DD",X"E5",X"FD",X"E5",X"D5",X"CD",X"A6",X"02",X"CD",X"66",X"03",X"CD",X"F8",X"03",X"CD",X"6D",
		X"04",X"CD",X"EE",X"04",X"3A",X"2F",X"F4",X"FE",X"09",X"38",X"05",X"3E",X"09",X"32",X"2F",X"F4",
		X"DB",X"00",X"E6",X"20",X"20",X"35",X"21",X"1E",X"F4",X"36",X"02",X"23",X"36",X"09",X"23",X"22",
		X"1B",X"F4",X"3E",X"02",X"32",X"1D",X"F4",X"CD",X"31",X"06",X"21",X"00",X"60",X"2B",X"7C",X"B5",
		X"20",X"FB",X"DB",X"00",X"E6",X"20",X"28",X"F2",X"3A",X"03",X"F0",X"E6",X"80",X"28",X"0A",X"3A",
		X"2F",X"F4",X"B7",X"28",X"04",X"3D",X"32",X"2F",X"F4",X"18",X"FE",X"D1",X"FD",X"E1",X"DD",X"E1",
		X"C1",X"E1",X"F1",X"FB",X"ED",X"4D",X"3A",X"A4",X"F0",X"F6",X"30",X"E6",X"B0",X"4F",X"D3",X"04",
		X"06",X"18",X"10",X"FE",X"DB",X"02",X"57",X"79",X"EE",X"80",X"4F",X"D3",X"04",X"06",X"20",X"10",
		X"FE",X"79",X"F6",X"70",X"32",X"A4",X"F0",X"D3",X"04",X"CB",X"79",X"28",X"21",X"06",X"05",X"3A",
		X"15",X"F0",X"B7",X"28",X"02",X"06",X"06",X"7A",X"0E",X"00",X"18",X"01",X"0C",X"90",X"30",X"FC",
		X"79",X"21",X"38",X"F4",X"96",X"30",X"01",X"AF",X"E6",X"3F",X"32",X"7E",X"F0",X"C9",X"3A",X"01",
		X"F4",X"B7",X"C0",X"21",X"37",X"F4",X"7A",X"ED",X"44",X"96",X"32",X"A2",X"F0",X"CB",X"2F",X"CB",
		X"2F",X"CB",X"2F",X"47",X"3A",X"03",X"F0",X"E6",X"16",X"C0",X"3A",X"14",X"F0",X"B7",X"28",X"09",
		X"3A",X"82",X"F0",X"CB",X"3F",X"3C",X"4F",X"18",X"10",X"3A",X"15",X"F0",X"B7",X"28",X"30",X"0E",
		X"03",X"3A",X"03",X"F0",X"E6",X"40",X"28",X"01",X"0C",X"21",X"A3",X"F0",X"35",X"C0",X"3A",X"A1",
		X"F0",X"B8",X"28",X"16",X"CB",X"7F",X"20",X"0A",X"CB",X"78",X"20",X"03",X"B8",X"38",X"0A",X"3D",
		X"18",X"08",X"CB",X"78",X"28",X"03",X"B8",X"30",X"F6",X"3C",X"47",X"79",X"32",X"A3",X"F0",X"78",
		X"CB",X"78",X"28",X"02",X"ED",X"44",X"FE",X"09",X"38",X"02",X"3E",X"08",X"CB",X"78",X"28",X"02",
		X"ED",X"44",X"32",X"A1",X"F0",X"C9",X"3A",X"5C",X"F0",X"F6",X"FB",X"57",X"3A",X"A4",X"F0",X"5F",
		X"3A",X"12",X"F0",X"A2",X"57",X"3A",X"A5",X"F0",X"AA",X"CA",X"D5",X"03",X"4F",X"CB",X"41",X"28",
		X"08",X"06",X"01",X"3E",X"04",X"CB",X"42",X"18",X"2F",X"CB",X"49",X"28",X"08",X"06",X"02",X"3E",
		X"03",X"CB",X"4A",X"18",X"23",X"CB",X"51",X"28",X"08",X"06",X"04",X"3E",X"02",X"CB",X"52",X"18",
		X"17",X"CB",X"59",X"28",X"08",X"06",X"08",X"3E",X"00",X"CB",X"5A",X"18",X"0B",X"CB",X"79",X"CA",
		X"D5",X"03",X"06",X"80",X"3E",X"01",X"CB",X"7A",X"28",X"02",X"F6",X"08",X"B3",X"50",X"D3",X"04",
		X"06",X"24",X"10",X"FE",X"E6",X"DF",X"D3",X"04",X"4F",X"3A",X"A5",X"F0",X"AA",X"32",X"A5",X"F0",
		X"79",X"F6",X"20",X"D3",X"04",X"3A",X"A6",X"F0",X"57",X"E6",X"F0",X"C8",X"7A",X"E6",X"0F",X"57",
		X"B3",X"D3",X"04",X"06",X"14",X"10",X"FE",X"E6",X"EF",X"D3",X"04",X"06",X"08",X"10",X"FE",X"F6",
		X"10",X"D3",X"04",X"7A",X"32",X"A6",X"F0",X"C9",X"21",X"0E",X"F4",X"DB",X"00",X"E6",X"01",X"BE",
		X"28",X"03",X"77",X"18",X"38",X"21",X"13",X"F4",X"B7",X"20",X"03",X"77",X"18",X"2F",X"BE",X"28",
		X"2C",X"77",X"DB",X"00",X"E6",X"80",X"28",X"25",X"2A",X"22",X"F6",X"23",X"22",X"22",X"F6",X"21",
		X"0A",X"F4",X"34",X"21",X"17",X"F4",X"34",X"3A",X"30",X"F4",X"3C",X"21",X"2B",X"F4",X"BE",X"38",
		X"09",X"21",X"2F",X"F4",X"3A",X"2C",X"F4",X"86",X"77",X"AF",X"32",X"30",X"F4",X"3A",X"0C",X"F4",
		X"3D",X"FA",X"55",X"04",X"32",X"0C",X"F4",X"FE",X"10",X"C0",X"3A",X"12",X"F4",X"CB",X"87",X"D3",
		X"00",X"32",X"12",X"F4",X"C9",X"3A",X"0A",X"F4",X"3D",X"F8",X"32",X"0A",X"F4",X"3E",X"20",X"32",
		X"0C",X"F4",X"3A",X"12",X"F4",X"CB",X"C7",X"D3",X"00",X"32",X"12",X"F4",X"C9",X"21",X"0F",X"F4",
		X"DB",X"00",X"E6",X"02",X"BE",X"28",X"03",X"77",X"18",X"44",X"21",X"14",X"F4",X"B7",X"20",X"03",
		X"77",X"18",X"3B",X"BE",X"28",X"38",X"77",X"DB",X"00",X"E6",X"80",X"28",X"31",X"2A",X"24",X"F6",
		X"23",X"22",X"24",X"F6",X"DB",X"03",X"E6",X"04",X"20",X"06",X"21",X"0B",X"F4",X"34",X"18",X"04",
		X"21",X"0A",X"F4",X"34",X"21",X"17",X"F4",X"34",X"3A",X"31",X"F4",X"3C",X"21",X"2D",X"F4",X"BE",
		X"38",X"09",X"21",X"2F",X"F4",X"3A",X"2E",X"F4",X"86",X"77",X"AF",X"32",X"31",X"F4",X"3A",X"0D",
		X"F4",X"3D",X"FA",X"D6",X"04",X"32",X"0D",X"F4",X"FE",X"10",X"C0",X"3A",X"12",X"F4",X"CB",X"8F",
		X"D3",X"00",X"32",X"12",X"F4",X"C9",X"3A",X"0B",X"F4",X"3D",X"F8",X"32",X"0B",X"F4",X"3E",X"20",
		X"32",X"0D",X"F4",X"3A",X"12",X"F4",X"CB",X"CF",X"D3",X"00",X"32",X"12",X"F4",X"C9",X"21",X"10",
		X"F4",X"DB",X"00",X"E6",X"40",X"BE",X"28",X"02",X"77",X"C9",X"21",X"15",X"F4",X"B7",X"20",X"03",
		X"77",X"18",X"12",X"BE",X"28",X"0F",X"77",X"DB",X"00",X"E6",X"80",X"28",X"08",X"21",X"17",X"F4",
		X"34",X"21",X"2F",X"F4",X"34",X"C9",X"3A",X"AB",X"F0",X"B7",X"CA",X"A4",X"05",X"AF",X"32",X"AB",
		X"F0",X"32",X"A0",X"F0",X"3A",X"15",X"F0",X"B7",X"28",X"04",X"21",X"90",X"F3",X"34",X"2A",X"A7",
		X"F0",X"01",X"83",X"C9",X"78",X"BC",X"20",X"1E",X"79",X"BD",X"20",X"1A",X"3E",X"01",X"32",X"A3",
		X"F0",X"32",X"14",X"F0",X"21",X"10",X"EA",X"36",X"00",X"01",X"83",X"00",X"11",X"0F",X"EA",X"ED",
		X"B8",X"CD",X"DD",X"05",X"18",X"2D",X"3A",X"14",X"F0",X"B7",X"C4",X"FD",X"05",X"2A",X"3C",X"F0",
		X"3E",X"1F",X"85",X"30",X"01",X"24",X"6F",X"7E",X"FE",X"69",X"20",X"0A",X"3E",X"01",X"32",X"E5",
		X"F0",X"32",X"E6",X"F0",X"18",X"0D",X"3A",X"8E",X"F3",X"FE",X"08",X"3E",X"00",X"38",X"01",X"3C",
		X"32",X"E5",X"F0",X"2A",X"A7",X"F0",X"DD",X"21",X"20",X"FA",X"06",X"10",X"11",X"02",X"00",X"7E",
		X"B7",X"28",X"03",X"1B",X"DD",X"23",X"23",X"7E",X"DD",X"77",X"00",X"DD",X"77",X"40",X"DD",X"19",
		X"23",X"10",X"E9",X"C9",X"3A",X"AC",X"F0",X"3C",X"E6",X"1F",X"32",X"AC",X"F0",X"06",X"A9",X"CB",
		X"5F",X"28",X"02",X"06",X"69",X"E6",X"0F",X"CB",X"3F",X"CB",X"27",X"21",X"21",X"06",X"85",X"30",
		X"01",X"24",X"6F",X"7E",X"DD",X"21",X"20",X"FA",X"DD",X"77",X"0C",X"DD",X"77",X"4C",X"23",X"7E",
		X"DD",X"77",X"14",X"DD",X"77",X"54",X"DD",X"70",X"04",X"DD",X"70",X"44",X"C9",X"06",X"40",X"21",
		X"45",X"E8",X"7E",X"B7",X"28",X"13",X"FE",X"01",X"20",X"04",X"3E",X"76",X"18",X"0A",X"FE",X"3A",
		X"30",X"04",X"D6",X"23",X"18",X"02",X"C6",X"1B",X"77",X"23",X"10",X"E6",X"C9",X"AF",X"32",X"14",
		X"F0",X"06",X"40",X"21",X"45",X"E8",X"7E",X"B7",X"28",X"13",X"FE",X"76",X"20",X"04",X"3E",X"01",
		X"18",X"0A",X"FE",X"5C",X"38",X"04",X"D6",X"1B",X"18",X"02",X"C6",X"23",X"77",X"23",X"10",X"E6",
		X"C9",X"21",X"2B",X"A1",X"23",X"69",X"1B",X"6A",X"1A",X"2B",X"21",X"23",X"A1",X"1B",X"69",X"1A",
		X"6A",X"21",X"17",X"F4",X"7E",X"B7",X"28",X"16",X"35",X"21",X"1D",X"F4",X"ED",X"5B",X"1B",X"F4",
		X"3E",X"02",X"12",X"13",X"34",X"3E",X"0C",X"12",X"13",X"ED",X"53",X"1B",X"F4",X"34",X"3A",X"1D",
		X"F4",X"B7",X"28",X"6E",X"0E",X"1D",X"21",X"1E",X"F4",X"06",X"01",X"57",X"7E",X"CB",X"7F",X"28",
		X"25",X"78",X"FE",X"01",X"28",X"0D",X"FE",X"03",X"3E",X"00",X"28",X"03",X"ED",X"79",X"0C",X"ED",
		X"79",X"18",X"21",X"06",X"03",X"7E",X"ED",X"79",X"23",X"0C",X"10",X"F9",X"7A",X"D6",X"03",X"28",
		X"36",X"30",X"14",X"AF",X"18",X"31",X"ED",X"79",X"23",X"0C",X"78",X"BA",X"28",X"1C",X"3C",X"47",
		X"FE",X"04",X"20",X"C8",X"05",X"7A",X"90",X"32",X"1D",X"F4",X"11",X"1E",X"F4",X"47",X"7E",X"12",
		X"13",X"23",X"10",X"FA",X"ED",X"53",X"1B",X"F4",X"18",X"28",X"3E",X"03",X"92",X"28",X"08",X"16",
		X"00",X"ED",X"51",X"0C",X"3D",X"20",X"FA",X"21",X"1E",X"F4",X"22",X"1B",X"F4",X"32",X"1D",X"F4",
		X"18",X"10",X"3A",X"1A",X"F4",X"E6",X"40",X"C8",X"0E",X"1D",X"06",X"03",X"AF",X"ED",X"79",X"0C",
		X"10",X"FB",X"3A",X"19",X"F4",X"EE",X"80",X"32",X"19",X"F4",X"21",X"1A",X"F4",X"B6",X"D3",X"1C",
		X"36",X"00",X"C9",X"3A",X"7A",X"F3",X"FE",X"01",X"20",X"71",X"21",X"7C",X"F3",X"35",X"20",X"6B",
		X"3A",X"03",X"F0",X"E6",X"03",X"3A",X"7D",X"F3",X"28",X"02",X"C6",X"02",X"77",X"06",X"03",X"21",
		X"81",X"F3",X"35",X"F2",X"4B",X"07",X"36",X"09",X"2B",X"10",X"F7",X"06",X"03",X"21",X"6E",X"E8",
		X"36",X"00",X"23",X"10",X"FB",X"21",X"70",X"E8",X"06",X"07",X"0E",X"00",X"3A",X"84",X"F3",X"B7",
		X"28",X"16",X"36",X"01",X"2B",X"05",X"0C",X"FE",X"02",X"30",X"07",X"3A",X"85",X"F3",X"FE",X"08",
		X"38",X"06",X"34",X"36",X"01",X"2B",X"05",X"0C",X"AF",X"77",X"2B",X"10",X"FB",X"32",X"7A",X"F3",
		X"79",X"32",X"89",X"F3",X"B7",X"C8",X"0E",X"0B",X"C3",X"4E",X"3D",X"06",X"03",X"21",X"6E",X"E8",
		X"11",X"81",X"F3",X"1A",X"F6",X"30",X"77",X"23",X"1B",X"10",X"F8",X"3A",X"5D",X"F3",X"B7",X"C0",
		X"3A",X"16",X"F4",X"B7",X"C0",X"3A",X"28",X"F0",X"B7",X"28",X"13",X"3A",X"29",X"F0",X"B7",X"C0",
		X"3C",X"32",X"29",X"F0",X"11",X"37",X"B9",X"21",X"7A",X"E8",X"CD",X"18",X"3F",X"C9",X"3A",X"29",
		X"F0",X"B7",X"28",X"0F",X"AF",X"32",X"29",X"F0",X"06",X"09",X"21",X"7A",X"E8",X"36",X"00",X"2B",
		X"10",X"FB",X"C9",X"3A",X"14",X"F0",X"B7",X"0E",X"30",X"28",X"02",X"0E",X"0D",X"06",X"06",X"21",
		X"7A",X"E8",X"11",X"82",X"F3",X"1A",X"B7",X"28",X"01",X"81",X"77",X"2B",X"13",X"1A",X"81",X"BE",
		X"28",X"01",X"77",X"10",X"F6",X"C9",X"CD",X"3A",X"3D",X"CD",X"3A",X"3D",X"DD",X"21",X"23",X"0A",
		X"CD",X"76",X"09",X"F5",X"CD",X"16",X"05",X"21",X"00",X"F8",X"36",X"FE",X"3E",X"01",X"32",X"5D",
		X"F3",X"AF",X"32",X"01",X"F4",X"CD",X"4C",X"09",X"CD",X"67",X"09",X"F1",X"B7",X"28",X"12",X"DD",
		X"21",X"FA",X"07",X"CD",X"97",X"0A",X"3E",X"01",X"32",X"5D",X"F3",X"CD",X"CB",X"0A",X"F6",X"01",
		X"C9",X"CD",X"CB",X"0A",X"C0",X"CD",X"64",X"0C",X"AF",X"C9",X"04",X"08",X"D8",X"E8",X"F8",X"E8",
		X"0E",X"08",X"12",X"08",X"52",X"41",X"4D",X"20",X"45",X"52",X"52",X"4F",X"52",X"00",X"42",X"32",
		X"20",X"00",X"46",X"36",X"20",X"00",X"F3",X"CD",X"B6",X"07",X"F5",X"21",X"16",X"F4",X"CD",X"2E",
		X"3D",X"21",X"1E",X"F4",X"22",X"1B",X"F4",X"F1",X"FB",X"28",X"25",X"21",X"59",X"EA",X"11",X"C0",
		X"08",X"CD",X"18",X"3F",X"21",X"99",X"EA",X"11",X"D7",X"08",X"CD",X"18",X"3F",X"3E",X"01",X"32",
		X"5D",X"F3",X"CD",X"AB",X"A3",X"20",X"09",X"DB",X"00",X"E6",X"80",X"C0",X"D3",X"E0",X"18",X"ED",
		X"CD",X"02",X"09",X"CD",X"67",X"09",X"3E",X"01",X"32",X"5D",X"F3",X"CD",X"85",X"0B",X"F5",X"0E",
		X"02",X"CD",X"4E",X"3D",X"CD",X"F9",X"3C",X"0E",X"02",X"CD",X"4E",X"3D",X"CD",X"F9",X"3C",X"F1",
		X"28",X"20",X"21",X"59",X"EA",X"11",X"C0",X"08",X"CD",X"18",X"3F",X"21",X"99",X"EA",X"11",X"D7",
		X"08",X"CD",X"18",X"3F",X"CD",X"AB",X"A3",X"20",X"09",X"DB",X"00",X"E6",X"80",X"C0",X"D3",X"E0",
		X"18",X"F2",X"CD",X"67",X"09",X"21",X"18",X"E9",X"11",X"E3",X"08",X"CD",X"18",X"3F",X"21",X"36",
		X"E9",X"11",X"FA",X"08",X"CD",X"18",X"3F",X"11",X"FF",X"FF",X"CD",X"AB",X"A3",X"C0",X"DB",X"00",
		X"E6",X"80",X"C0",X"D3",X"E0",X"1B",X"7A",X"B3",X"20",X"F0",X"CD",X"67",X"09",X"C3",X"16",X"08",
		X"48",X"49",X"54",X"20",X"57",X"45",X"41",X"50",X"4F",X"4E",X"53",X"20",X"56",X"41",X"4E",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"54",X"4F",X"20",X"43",X"4F",X"4E",X"54",X"49",X"4E",
		X"55",X"45",X"00",X"48",X"49",X"54",X"20",X"57",X"45",X"41",X"50",X"4F",X"4E",X"53",X"20",X"56",
		X"41",X"4E",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"54",X"4F",X"20",X"45",X"58",X"49",
		X"54",X"00",X"CD",X"4C",X"09",X"CD",X"67",X"09",X"CD",X"F9",X"3C",X"06",X"0A",X"21",X"38",X"09",
		X"DD",X"21",X"20",X"FA",X"7E",X"B7",X"28",X"02",X"DD",X"23",X"23",X"7E",X"DD",X"77",X"00",X"CD",
		X"2C",X"09",X"DD",X"77",X"40",X"CD",X"2C",X"09",X"23",X"10",X"E5",X"C9",X"F5",X"C5",X"06",X"14",
		X"CD",X"F9",X"3C",X"10",X"FB",X"C1",X"F1",X"C9",X"00",X"20",X"00",X"7C",X"00",X"05",X"01",X"C7",
		X"01",X"D0",X"01",X"30",X"01",X"E8",X"01",X"FF",X"00",X"00",X"00",X"00",X"DD",X"21",X"20",X"FA",
		X"DD",X"36",X"00",X"49",X"DD",X"36",X"40",X"49",X"21",X"00",X"E0",X"01",X"FF",X"07",X"36",X"04",
		X"23",X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"21",X"00",X"E8",X"01",X"FF",X"03",X"36",X"00",X"23",
		X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"AF",X"F5",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"7C",X"B5",
		X"20",X"02",X"F1",X"C9",X"DD",X"5E",X"04",X"DD",X"56",X"05",X"DD",X"4E",X"02",X"DD",X"46",X"03",
		X"ED",X"B0",X"DD",X"7E",X"07",X"32",X"FF",X"F7",X"D3",X"E0",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",X"B3",X"28",X"11",X"06",X"02",X"3E",X"00",X"77",X"BE",
		X"C2",X"1E",X"0A",X"F6",X"FF",X"10",X"F7",X"23",X"1B",X"18",X"EB",X"DD",X"66",X"01",X"DD",X"6E",
		X"00",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"D3",X"E0",X"7A",X"B3",X"28",X"06",X"36",X"00",X"23",
		X"1B",X"18",X"F6",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"7A",
		X"B3",X"28",X"15",X"7E",X"FE",X"00",X"C2",X"1E",X"0A",X"3E",X"01",X"77",X"BE",X"C2",X"1E",X"0A",
		X"CB",X"27",X"30",X"F7",X"23",X"1B",X"18",X"E7",X"AF",X"DD",X"66",X"05",X"DD",X"6E",X"04",X"DD",
		X"56",X"01",X"DD",X"5E",X"00",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"D3",X"E0",X"ED",X"B0",X"47",
		X"F1",X"AF",X"32",X"FF",X"F7",X"B0",X"11",X"08",X"00",X"DD",X"19",X"C3",X"77",X"09",X"DD",X"7E",
		X"06",X"18",X"D6",X"00",X"F0",X"00",X"02",X"00",X"F2",X"01",X"01",X"00",X"F2",X"00",X"02",X"00",
		X"F0",X"01",X"02",X"00",X"F4",X"00",X"02",X"00",X"F2",X"01",X"03",X"00",X"F6",X"FF",X"01",X"00",
		X"F0",X"01",X"04",X"00",X"E0",X"00",X"04",X"00",X"F0",X"20",X"05",X"00",X"E4",X"00",X"04",X"00",
		X"F0",X"20",X"05",X"00",X"E8",X"00",X"04",X"00",X"F0",X"20",X"06",X"00",X"00",X"3A",X"FF",X"F7",
		X"B7",X"C8",X"DD",X"21",X"23",X"0A",X"11",X"08",X"00",X"47",X"DD",X"7E",X"07",X"B8",X"28",X"0C",
		X"DD",X"19",X"DD",X"7E",X"00",X"DD",X"B6",X"01",X"20",X"F0",X"18",X"17",X"DD",X"66",X"05",X"DD",
		X"6E",X"04",X"DD",X"56",X"01",X"DD",X"5E",X"00",X"DD",X"4E",X"02",X"DD",X"46",X"03",X"D3",X"E0",
		X"ED",X"B0",X"AF",X"32",X"FF",X"F7",X"C9",X"F5",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"5E",
		X"00",X"DD",X"56",X"01",X"CD",X"18",X"3F",X"F1",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"01",X"06",
		X"00",X"DD",X"09",X"CB",X"3F",X"30",X"0B",X"DD",X"5E",X"00",X"DD",X"56",X"01",X"F5",X"CD",X"18",
		X"3F",X"F1",X"01",X"02",X"00",X"DD",X"09",X"B7",X"20",X"E9",X"C9",X"3E",X"01",X"32",X"5D",X"F3",
		X"DD",X"21",X"0F",X"0B",X"16",X"00",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"DD",X"4E",X"00",X"DD",
		X"46",X"01",X"78",X"B1",X"28",X"1C",X"AF",X"86",X"23",X"0D",X"20",X"FB",X"05",X"20",X"F8",X"DD",
		X"BE",X"04",X"28",X"05",X"7A",X"DD",X"B6",X"05",X"57",X"01",X"06",X"00",X"DD",X"09",X"D3",X"E0",
		X"18",X"D4",X"7A",X"B7",X"C8",X"DD",X"21",X"36",X"0B",X"CD",X"97",X"0A",X"F6",X"01",X"C9",X"00",
		X"20",X"00",X"00",X"81",X"01",X"00",X"20",X"00",X"20",X"05",X"02",X"00",X"20",X"00",X"40",X"74",
		X"04",X"00",X"20",X"00",X"60",X"95",X"08",X"00",X"20",X"00",X"80",X"A0",X"10",X"00",X"40",X"00",
		X"A0",X"93",X"20",X"00",X"00",X"7F",X"4A",X"0B",X"36",X"E9",X"55",X"E9",X"54",X"0B",X"58",X"0B",
		X"5C",X"0B",X"60",X"0B",X"64",X"0B",X"68",X"0B",X"6C",X"0B",X"52",X"4F",X"4D",X"20",X"45",X"52",
		X"52",X"4F",X"52",X"00",X"44",X"32",X"20",X"00",X"44",X"33",X"20",X"00",X"44",X"34",X"20",X"00",
		X"44",X"35",X"20",X"00",X"44",X"36",X"20",X"00",X"44",X"37",X"20",X"00",X"44",X"38",X"20",X"00",
		X"CD",X"3A",X"3D",X"CD",X"64",X"0C",X"CD",X"F9",X"3C",X"DB",X"00",X"E6",X"80",X"20",X"05",X"CD",
		X"AB",X"A3",X"28",X"F2",X"C9",X"0E",X"02",X"CD",X"4E",X"3D",X"CD",X"F9",X"3C",X"CD",X"F9",X"3C",
		X"CD",X"F9",X"3C",X"CD",X"67",X"09",X"CD",X"3A",X"3D",X"0E",X"02",X"CD",X"4E",X"3D",X"0E",X"06",
		X"CD",X"4E",X"3D",X"CD",X"F9",X"3C",X"CD",X"F9",X"3C",X"DD",X"21",X"12",X"0C",X"01",X"00",X"04",
		X"CD",X"F9",X"3C",X"C5",X"0E",X"1F",X"DD",X"7E",X"00",X"06",X"04",X"ED",X"79",X"0D",X"10",X"FB",
		X"CD",X"F9",X"3C",X"CD",X"F9",X"3C",X"DB",X"07",X"C1",X"DD",X"BE",X"00",X"28",X"01",X"0C",X"DD",
		X"23",X"10",X"E0",X"79",X"B7",X"28",X"05",X"11",X"16",X"0C",X"18",X"10",X"06",X"64",X"DB",X"07",
		X"E6",X"80",X"28",X"19",X"CD",X"F9",X"3C",X"10",X"F5",X"11",X"26",X"0C",X"21",X"D9",X"EA",X"CD",
		X"18",X"3F",X"21",X"B9",X"EA",X"11",X"34",X"0C",X"CD",X"18",X"3F",X"18",X"0B",X"DB",X"07",X"B7",
		X"C8",X"DD",X"21",X"40",X"0C",X"CD",X"97",X"0A",X"06",X"60",X"CD",X"F9",X"3C",X"10",X"FB",X"F6",
		X"01",X"C9",X"00",X"FF",X"55",X"AA",X"49",X"4E",X"54",X"45",X"52",X"46",X"41",X"43",X"45",X"20",
		X"45",X"52",X"52",X"4F",X"52",X"00",X"42",X"4F",X"41",X"52",X"44",X"20",X"54",X"49",X"4D",X"45",
		X"4F",X"55",X"54",X"00",X"53",X"4F",X"55",X"4E",X"44",X"20",X"42",X"4F",X"41",X"52",X"44",X"00",
		X"34",X"0C",X"B9",X"EA",X"D9",X"EA",X"50",X"0C",X"54",X"0C",X"58",X"0C",X"5C",X"0C",X"61",X"0C",
		X"41",X"37",X"20",X"00",X"41",X"38",X"20",X"00",X"41",X"39",X"20",X"00",X"41",X"31",X"30",X"20",
		X"00",X"41",X"36",X"00",X"CD",X"4C",X"09",X"21",X"00",X"E8",X"01",X"FF",X"03",X"36",X"23",X"23",
		X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"3A",X"0A",X"F0",X"B7",X"C0",X"3A",X"15",X"F0",X"21",X"16",
		X"F0",X"BE",X"C0",X"3A",X"06",X"F0",X"FE",X"02",X"D2",X"0F",X"0D",X"21",X"57",X"F0",X"7E",X"FE",
		X"01",X"38",X"7C",X"28",X"03",X"35",X"18",X"77",X"3A",X"60",X"F0",X"B7",X"28",X"1A",X"DD",X"E5",
		X"DD",X"2A",X"5F",X"F0",X"DD",X"7E",X"02",X"FE",X"06",X"38",X"0A",X"DD",X"7E",X"01",X"B7",X"28",
		X"04",X"DD",X"E1",X"18",X"5A",X"DD",X"E1",X"AF",X"32",X"57",X"F0",X"21",X"33",X"F0",X"7E",X"FE",
		X"04",X"38",X"02",X"36",X"03",X"32",X"34",X"F0",X"DD",X"22",X"5F",X"F0",X"DD",X"36",X"06",X"29",
		X"3E",X"06",X"32",X"59",X"F0",X"3A",X"5B",X"F0",X"B7",X"28",X"0E",X"DD",X"36",X"01",X"81",X"DD",
		X"36",X"03",X"00",X"DD",X"36",X"0B",X"00",X"18",X"10",X"DD",X"36",X"01",X"80",X"3A",X"82",X"F0",
		X"C6",X"03",X"DD",X"77",X"03",X"DD",X"36",X"0B",X"0E",X"3E",X"1F",X"2A",X"3C",X"F0",X"85",X"30",
		X"01",X"24",X"6F",X"7E",X"DD",X"77",X"1D",X"2B",X"7E",X"DD",X"77",X"02",X"C3",X"F5",X"0D",X"21",
		X"45",X"F0",X"7E",X"FE",X"01",X"38",X"33",X"28",X"03",X"35",X"18",X"2E",X"3A",X"82",X"F0",X"FE",
		X"0F",X"30",X"27",X"FE",X"05",X"38",X"23",X"3A",X"49",X"F0",X"B7",X"20",X"1D",X"36",X"00",X"3A",
		X"15",X"F0",X"B7",X"28",X"08",X"3A",X"90",X"F3",X"B7",X"28",X"0F",X"18",X"05",X"3E",X"01",X"32",
		X"46",X"F0",X"DD",X"22",X"48",X"F0",X"3E",X"09",X"18",X"3A",X"3A",X"01",X"F4",X"06",X"07",X"B7",
		X"28",X"02",X"06",X"03",X"CD",X"E7",X"3C",X"A0",X"47",X"3A",X"15",X"F0",X"B7",X"20",X"23",X"3A",
		X"8E",X"F3",X"FE",X"05",X"38",X"1C",X"D6",X"02",X"B8",X"38",X"17",X"78",X"E6",X"03",X"47",X"3A",
		X"14",X"F0",X"B7",X"3E",X"08",X"20",X"02",X"3E",X"0A",X"80",X"32",X"37",X"F0",X"78",X"E6",X"01",
		X"18",X"02",X"04",X"78",X"47",X"CB",X"27",X"80",X"C6",X"02",X"2A",X"3C",X"F0",X"85",X"30",X"01",
		X"24",X"6F",X"7E",X"B7",X"20",X"11",X"3A",X"15",X"F0",X"21",X"FA",X"B9",X"28",X"03",X"21",X"C0",
		X"BA",X"22",X"3C",X"F0",X"AF",X"18",X"B1",X"DD",X"77",X"06",X"3C",X"DD",X"77",X"1D",X"2B",X"7E",
		X"B7",X"20",X"2C",X"3A",X"15",X"F0",X"B7",X"20",X"14",X"3A",X"42",X"F0",X"B7",X"28",X"0E",X"DD",
		X"36",X"01",X"81",X"DD",X"36",X"03",X"00",X"DD",X"36",X"0B",X"00",X"18",X"23",X"DD",X"36",X"01",
		X"80",X"3A",X"82",X"F0",X"C6",X"02",X"DD",X"77",X"03",X"DD",X"36",X"0B",X"0E",X"18",X"11",X"FE",
		X"FF",X"38",X"03",X"3A",X"37",X"F0",X"DD",X"77",X"0B",X"DD",X"77",X"03",X"DD",X"36",X"01",X"80",
		X"2B",X"7E",X"DD",X"77",X"02",X"E6",X"0F",X"47",X"21",X"E1",X"BA",X"85",X"30",X"01",X"24",X"6F",
		X"7E",X"DD",X"77",X"0E",X"21",X"EA",X"BA",X"78",X"85",X"30",X"01",X"24",X"6F",X"7E",X"DD",X"77",
		X"0F",X"DD",X"36",X"0D",X"01",X"DD",X"36",X"0C",X"01",X"DD",X"36",X"04",X"00",X"3E",X"20",X"DD",
		X"77",X"11",X"3A",X"82",X"F0",X"DD",X"BE",X"03",X"30",X"0A",X"DD",X"36",X"08",X"01",X"DD",X"36",
		X"07",X"20",X"18",X"0E",X"3A",X"9F",X"F0",X"B7",X"20",X"F0",X"DD",X"36",X"08",X"FF",X"DD",X"36",
		X"07",X"E0",X"06",X"00",X"DD",X"70",X"05",X"DD",X"70",X"0A",X"DD",X"70",X"1F",X"DD",X"70",X"1C",
		X"DD",X"70",X"1E",X"DD",X"70",X"21",X"DD",X"36",X"22",X"01",X"DD",X"7E",X"13",X"B7",X"28",X"08",
		X"DD",X"70",X"13",X"67",X"DD",X"6E",X"12",X"70",X"DD",X"7E",X"15",X"B7",X"28",X"08",X"DD",X"70",
		X"15",X"67",X"DD",X"6E",X"14",X"70",X"DD",X"7E",X"18",X"B7",X"28",X"08",X"DD",X"70",X"18",X"67",
		X"DD",X"6E",X"17",X"70",X"DD",X"7E",X"09",X"FE",X"03",X"20",X"08",X"21",X"F4",X"F8",X"70",X"21",
		X"F8",X"F8",X"70",X"DD",X"36",X"09",X"FF",X"21",X"32",X"F0",X"34",X"C9",X"21",X"82",X"F0",X"DD",
		X"7E",X"01",X"E6",X"0F",X"C2",X"DD",X"0F",X"DD",X"35",X"0D",X"C2",X"DD",X"0F",X"DD",X"7E",X"02",
		X"47",X"E6",X"0F",X"C2",X"4D",X"0F",X"CB",X"78",X"28",X"25",X"DD",X"7E",X"08",X"B7",X"C2",X"48",
		X"0F",X"3A",X"01",X"F0",X"D6",X"40",X"DD",X"BE",X"07",X"DD",X"46",X"0B",X"7E",X"30",X"02",X"C6",
		X"02",X"B8",X"38",X"01",X"78",X"DD",X"77",X"03",X"DD",X"36",X"0D",X"01",X"C3",X"DD",X"0F",X"3A",
		X"46",X"F0",X"B7",X"CA",X"B1",X"0F",X"CD",X"E7",X"3C",X"E5",X"21",X"47",X"F0",X"A6",X"3C",X"DD",
		X"77",X"0D",X"E1",X"3A",X"03",X"F0",X"E6",X"13",X"C2",X"DD",X"0F",X"DD",X"7E",X"08",X"B7",X"20",
		X"47",X"3A",X"00",X"F0",X"DD",X"96",X"05",X"30",X"02",X"ED",X"44",X"FE",X"14",X"30",X"0A",X"DD",
		X"7E",X"07",X"FE",X"E0",X"30",X"03",X"7E",X"18",X"1D",X"3A",X"01",X"F0",X"D6",X"0A",X"DD",X"BE",
		X"07",X"CA",X"DD",X"0F",X"7E",X"38",X"0B",X"FE",X"02",X"38",X"01",X"3D",X"DD",X"77",X"03",X"C3",
		X"DD",X"0F",X"DD",X"7E",X"03",X"3C",X"DD",X"BE",X"0B",X"38",X"03",X"DD",X"7E",X"0B",X"DD",X"77",
		X"03",X"DD",X"36",X"0D",X"04",X"C3",X"DD",X"0F",X"CB",X"27",X"86",X"18",X"E9",X"FE",X"06",X"38",
		X"60",X"DD",X"36",X"0D",X"01",X"DD",X"7E",X"09",X"FE",X"FF",X"28",X"11",X"3A",X"06",X"F0",X"DD",
		X"BE",X"09",X"C2",X"DD",X"0F",X"3A",X"03",X"F0",X"E6",X"03",X"C2",X"DD",X"0F",X"DD",X"7E",X"08",
		X"B7",X"28",X"15",X"CB",X"27",X"CB",X"27",X"86",X"CB",X"7F",X"28",X"07",X"3E",X"02",X"32",X"5B",
		X"F0",X"3E",X"0A",X"DD",X"77",X"03",X"18",X"55",X"3A",X"00",X"F0",X"DD",X"96",X"05",X"30",X"02",
		X"ED",X"44",X"FE",X"14",X"30",X"0A",X"DD",X"7E",X"07",X"FE",X"E0",X"30",X"03",X"7E",X"18",X"96",
		X"3A",X"01",X"F0",X"D6",X"38",X"DD",X"BE",X"07",X"38",X"88",X"7E",X"B7",X"20",X"88",X"3C",X"18",
		X"85",X"CD",X"E7",X"3C",X"E6",X"1F",X"3C",X"DD",X"77",X"0D",X"E6",X"01",X"47",X"DD",X"7E",X"0B",
		X"DD",X"BE",X"03",X"28",X"0B",X"38",X"0F",X"DD",X"34",X"03",X"DD",X"36",X"0D",X"02",X"18",X"0D",
		X"90",X"DD",X"77",X"03",X"18",X"07",X"DD",X"35",X"03",X"DD",X"36",X"0D",X"02",X"DD",X"7E",X"08",
		X"47",X"3A",X"D8",X"F0",X"B7",X"28",X"1C",X"78",X"FE",X"01",X"28",X"0C",X"30",X"15",X"DD",X"7E",
		X"05",X"B7",X"20",X"0F",X"06",X"01",X"18",X"07",X"DD",X"7E",X"07",X"FE",X"80",X"30",X"04",X"DD",
		X"36",X"07",X"80",X"7E",X"DD",X"96",X"03",X"DD",X"77",X"10",X"30",X"08",X"DD",X"86",X"07",X"38",
		X"6F",X"05",X"18",X"6C",X"20",X"64",X"7E",X"B7",X"20",X"30",X"DD",X"7E",X"01",X"E6",X"0A",X"20",
		X"58",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"06",X"38",X"10",X"3A",X"58",X"F0",X"FE",X"05",X"30",
		X"48",X"3E",X"01",X"2F",X"DD",X"A6",X"01",X"DD",X"77",X"01",X"DD",X"36",X"03",X"05",X"DD",X"7E",
		X"04",X"B7",X"20",X"BF",X"DD",X"36",X"04",X"02",X"18",X"B9",X"DD",X"7E",X"01",X"E6",X"0A",X"20",
		X"28",X"DD",X"7E",X"02",X"E6",X"0F",X"28",X"21",X"FE",X"05",X"30",X"1D",X"78",X"FE",X"01",X"38",
		X"18",X"DD",X"7E",X"03",X"28",X"08",X"D6",X"02",X"30",X"06",X"7E",X"3C",X"18",X"02",X"C6",X"02",
		X"DD",X"77",X"03",X"DD",X"36",X"0D",X"02",X"18",X"8A",X"AF",X"DD",X"86",X"07",X"30",X"01",X"04",
		X"4F",X"78",X"FE",X"01",X"DA",X"94",X"11",X"28",X"22",X"DD",X"7E",X"02",X"E6",X"10",X"79",X"20",
		X"07",X"FE",X"F8",X"D2",X"A7",X"11",X"18",X"05",X"FE",X"E8",X"D2",X"A7",X"11",X"DD",X"7E",X"05",
		X"B7",X"20",X"0E",X"79",X"FE",X"40",X"38",X"75",X"C3",X"A0",X"11",X"DD",X"7E",X"05",X"B7",X"28",
		X"66",X"DD",X"77",X"0A",X"DD",X"36",X"05",X"00",X"DD",X"7E",X"18",X"B7",X"28",X"0A",X"67",X"DD",
		X"6E",X"17",X"36",X"00",X"DD",X"36",X"18",X"00",X"DD",X"7E",X"13",X"B7",X"28",X"0A",X"67",X"DD",
		X"6E",X"12",X"36",X"00",X"DD",X"36",X"13",X"00",X"DD",X"7E",X"15",X"B7",X"28",X"0A",X"67",X"DD",
		X"6E",X"14",X"36",X"00",X"DD",X"36",X"15",X"00",X"DD",X"7E",X"01",X"E6",X"04",X"28",X"0F",X"DD",
		X"7E",X"0C",X"FE",X"14",X"38",X"08",X"DD",X"7E",X"02",X"CD",X"91",X"3E",X"18",X"1F",X"DD",X"7E",
		X"02",X"E6",X"0F",X"20",X"08",X"3A",X"06",X"F0",X"DD",X"BE",X"09",X"20",X"10",X"DD",X"7E",X"01",
		X"E6",X"0A",X"20",X"09",X"C3",X"A0",X"11",X"79",X"FE",X"C1",X"DA",X"A0",X"11",X"DD",X"7E",X"02",
		X"E6",X"0F",X"20",X"27",X"32",X"49",X"F0",X"32",X"46",X"F0",X"CD",X"01",X"56",X"3A",X"42",X"F0",
		X"B7",X"28",X"58",X"AF",X"32",X"42",X"F0",X"DD",X"7E",X"01",X"E6",X"02",X"20",X"4D",X"DD",X"7E",
		X"03",X"B7",X"20",X"47",X"21",X"45",X"F0",X"36",X"05",X"18",X"40",X"FE",X"06",X"38",X"3C",X"AF",
		X"32",X"58",X"F0",X"32",X"60",X"F0",X"3A",X"33",X"F0",X"FE",X"03",X"20",X"06",X"3A",X"34",X"F0",
		X"32",X"33",X"F0",X"21",X"5B",X"F0",X"7E",X"B7",X"28",X"13",X"47",X"DD",X"7E",X"01",X"E6",X"02",
		X"20",X"09",X"05",X"70",X"21",X"57",X"F0",X"36",X"03",X"18",X"10",X"36",X"00",X"3A",X"5E",X"F0",
		X"B7",X"28",X"05",X"3A",X"12",X"F0",X"E6",X"04",X"32",X"5C",X"F0",X"DD",X"36",X"01",X"00",X"21",
		X"32",X"F0",X"35",X"C9",X"79",X"FE",X"F8",X"38",X"0E",X"DD",X"7E",X"05",X"B7",X"C2",X"B1",X"10",
		X"DD",X"70",X"08",X"DD",X"71",X"07",X"C9",X"DD",X"7E",X"05",X"B7",X"3E",X"10",X"28",X"08",X"DD",
		X"70",X"08",X"DD",X"71",X"07",X"3E",X"20",X"DD",X"B6",X"01",X"DD",X"77",X"01",X"C9",X"21",X"BE",
		X"06",X"22",X"91",X"F0",X"7D",X"D3",X"84",X"7C",X"D3",X"85",X"AF",X"D3",X"86",X"DD",X"21",X"00",
		X"F8",X"DD",X"36",X"00",X"FE",X"DD",X"77",X"01",X"DD",X"77",X"02",X"DD",X"77",X"03",X"3E",X"8F",
		X"32",X"A5",X"F0",X"3E",X"02",X"32",X"7C",X"F3",X"32",X"7A",X"F3",X"DB",X"03",X"E6",X"01",X"3E",
		X"03",X"20",X"01",X"3D",X"32",X"7D",X"F3",X"21",X"04",X"F0",X"36",X"14",X"21",X"05",X"F0",X"36",
		X"04",X"21",X"07",X"F0",X"36",X"D3",X"21",X"06",X"F0",X"36",X"02",X"21",X"03",X"F0",X"36",X"80",
		X"21",X"13",X"F0",X"36",X"01",X"AF",X"32",X"11",X"F0",X"DD",X"21",X"74",X"F8",X"DD",X"36",X"02",
		X"0E",X"06",X"30",X"11",X"04",X"00",X"DD",X"21",X"FC",X"F8",X"DD",X"19",X"DD",X"36",X"02",X"19",
		X"10",X"F8",X"06",X"00",X"21",X"82",X"F2",X"70",X"2B",X"70",X"2B",X"70",X"2B",X"3A",X"34",X"F4",
		X"77",X"2B",X"3A",X"33",X"F4",X"77",X"2B",X"70",X"2B",X"70",X"21",X"89",X"F2",X"70",X"2B",X"70",
		X"2B",X"70",X"2B",X"3A",X"36",X"F4",X"77",X"2B",X"3A",X"35",X"F4",X"77",X"2B",X"70",X"2B",X"70",
		X"21",X"8A",X"F2",X"36",X"04",X"AF",X"32",X"49",X"F0",X"21",X"F3",X"BA",X"3A",X"32",X"F4",X"3D",
		X"CB",X"27",X"85",X"30",X"01",X"24",X"6F",X"5E",X"23",X"56",X"ED",X"53",X"30",X"F0",X"1A",X"32",
		X"33",X"F0",X"21",X"39",X"F0",X"36",X"0E",X"21",X"47",X"F0",X"36",X"1F",X"21",X"4D",X"F0",X"36",
		X"04",X"21",X"FC",X"F0",X"36",X"04",X"21",X"DD",X"F0",X"36",X"20",X"21",X"40",X"F0",X"36",X"04",
		X"11",X"03",X"00",X"AF",X"DD",X"21",X"61",X"F0",X"DD",X"77",X"00",X"DD",X"19",X"3C",X"FE",X"09",
		X"20",X"F6",X"DD",X"21",X"47",X"BC",X"DD",X"22",X"99",X"F0",X"DD",X"6E",X"00",X"DD",X"66",X"01",
		X"22",X"A7",X"F0",X"21",X"AB",X"F0",X"36",X"01",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"22",X"3C",
		X"F0",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"5E",X"23",X"56",X"ED",X"53",X"95",X"F0",X"23",X"7E",
		X"DD",X"21",X"61",X"F0",X"DD",X"77",X"01",X"DD",X"36",X"02",X"40",X"01",X"03",X"00",X"ED",X"43",
		X"7C",X"F0",X"23",X"23",X"E5",X"DD",X"E1",X"21",X"FE",X"03",X"22",X"97",X"F0",X"06",X"80",X"CD",
		X"41",X"46",X"10",X"FB",X"DD",X"22",X"93",X"F0",X"3E",X"00",X"DD",X"21",X"8B",X"F2",X"11",X"23",
		X"00",X"DD",X"77",X"00",X"DD",X"36",X"01",X"00",X"DD",X"19",X"3C",X"FE",X"06",X"20",X"F2",X"3A",
		X"35",X"F0",X"32",X"36",X"F0",X"C9",X"21",X"2B",X"F4",X"06",X"04",X"7E",X"B7",X"28",X"66",X"FE",
		X"0A",X"30",X"62",X"23",X"10",X"F5",X"7E",X"23",X"FE",X"0A",X"30",X"59",X"3A",X"2B",X"F4",X"BE",
		X"38",X"53",X"28",X"51",X"23",X"3A",X"2D",X"F4",X"BE",X"38",X"4A",X"28",X"48",X"23",X"23",X"23",
		X"23",X"23",X"23",X"23",X"23",X"06",X"07",X"7E",X"FE",X"0A",X"30",X"39",X"23",X"10",X"F8",X"06",
		X"1E",X"0E",X"03",X"7E",X"0D",X"20",X"04",X"0E",X"03",X"18",X"0C",X"FE",X"20",X"28",X"08",X"FE",
		X"41",X"38",X"22",X"FE",X"5B",X"30",X"1E",X"23",X"10",X"E9",X"01",X"98",X"01",X"21",X"62",X"F4",
		X"7E",X"E6",X"F0",X"FE",X"A0",X"30",X"0E",X"7E",X"E6",X"0F",X"FE",X"0A",X"30",X"07",X"23",X"0B",
		X"78",X"B1",X"20",X"EC",X"C9",X"11",X"2B",X"F4",X"21",X"BC",X"13",X"01",X"67",X"00",X"ED",X"B0",
		X"DB",X"03",X"E6",X"08",X"20",X"09",X"21",X"2B",X"F4",X"36",X"01",X"23",X"23",X"36",X"01",X"AF",
		X"01",X"94",X"01",X"AF",X"12",X"13",X"0B",X"78",X"B1",X"20",X"F8",X"C9",X"02",X"01",X"02",X"01",
		X"00",X"00",X"00",X"03",X"03",X"00",X"03",X"00",X"8C",X"0B",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"54",X"46",X"4C",X"4B",X"4F",X"20",X"47",X"47",X"20",X"41",X"47",X"20",X"52",X"4D",X"4C",
		X"53",X"50",X"20",X"53",X"56",X"20",X"42",X"46",X"43",X"4A",X"43",X"4B",X"53",X"4A",X"55",X"00",
		X"01",X"09",X"00",X"01",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"01",X"90",X"00",X"00",X"01",X"80",X"00",X"00",X"01",X"70",X"00",X"00",X"01",X"60",X"00",X"00",
		X"01",X"50",X"00",X"00",X"01",X"40",X"00",X"00",X"01",X"30",X"00",X"00",X"01",X"20",X"00",X"00",
		X"01",X"10",X"00",X"D5",X"DD",X"7E",X"01",X"EE",X"20",X"DD",X"77",X"01",X"47",X"3A",X"0A",X"F0",
		X"B7",X"28",X"09",X"3A",X"0C",X"F0",X"DD",X"86",X"05",X"C3",X"1B",X"1B",X"78",X"E6",X"0C",X"C2",
		X"30",X"19",X"78",X"E6",X"02",X"C2",X"0F",X"1B",X"DD",X"7E",X"03",X"B7",X"CA",X"B7",X"1B",X"3A",
		X"D8",X"F0",X"B7",X"28",X"35",X"DD",X"7E",X"08",X"B7",X"20",X"2F",X"3A",X"06",X"F0",X"DD",X"BE",
		X"09",X"20",X"27",X"3A",X"01",X"F0",X"C6",X"18",X"DD",X"BE",X"07",X"30",X"1D",X"3A",X"82",X"F0",
		X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"03",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"06",X"3E",X"80",
		X"38",X"02",X"3E",X"04",X"DD",X"77",X"0D",X"C3",X"0F",X"1B",X"CD",X"F3",X"43",X"DD",X"7E",X"05",
		X"DD",X"86",X"04",X"47",X"FD",X"21",X"5B",X"F2",X"CD",X"62",X"45",X"DA",X"21",X"15",X"DD",X"7E",
		X"02",X"E6",X"0F",X"FE",X"06",X"38",X"14",X"3A",X"58",X"F0",X"FE",X"05",X"38",X"0D",X"79",X"B7",
		X"28",X"09",X"DD",X"36",X"0D",X"01",X"DD",X"35",X"03",X"18",X"69",X"3A",X"06",X"F0",X"DD",X"BE",
		X"09",X"28",X"1B",X"3A",X"15",X"F0",X"B7",X"20",X"15",X"3A",X"55",X"F0",X"CB",X"5F",X"20",X"0E",
		X"E6",X"0F",X"FE",X"06",X"38",X"08",X"3E",X"02",X"20",X"01",X"2F",X"C3",X"EE",X"1A",X"DD",X"7E",
		X"0D",X"FE",X"04",X"30",X"04",X"DD",X"36",X"0D",X"04",X"DD",X"7E",X"0B",X"D6",X"03",X"DD",X"BE",
		X"03",X"30",X"03",X"DD",X"77",X"03",X"DD",X"36",X"0C",X"04",X"16",X"02",X"3A",X"15",X"F0",X"B7",
		X"28",X"0E",X"DD",X"7E",X"10",X"CB",X"7F",X"28",X"02",X"ED",X"44",X"B7",X"20",X"01",X"3C",X"57",
		X"79",X"B7",X"7A",X"0E",X"20",X"28",X"04",X"ED",X"44",X"0E",X"E0",X"DD",X"71",X"11",X"C3",X"EE",
		X"1A",X"DD",X"71",X"09",X"16",X"FF",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"06",X"38",X"08",X"3A",
		X"58",X"F0",X"FE",X"05",X"D2",X"15",X"16",X"1E",X"00",X"FD",X"21",X"8B",X"F2",X"7B",X"FE",X"06",
		X"CA",X"15",X"16",X"FD",X"7E",X"00",X"DD",X"BE",X"00",X"CA",X"0C",X"16",X"FD",X"7E",X"05",X"B7",
		X"CA",X"0C",X"16",X"DD",X"7E",X"10",X"FD",X"96",X"10",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"47",
		X"DD",X"7E",X"08",X"B7",X"20",X"3A",X"FD",X"B6",X"08",X"20",X"23",X"DD",X"7E",X"07",X"DD",X"86",
		X"0E",X"38",X"06",X"FD",X"BE",X"07",X"DA",X"0C",X"16",X"78",X"ED",X"44",X"FD",X"86",X"0E",X"C6",
		X"10",X"FD",X"86",X"07",X"38",X"2E",X"DD",X"BE",X"07",X"DA",X"0C",X"16",X"18",X"26",X"78",X"ED",
		X"44",X"FD",X"86",X"0E",X"C6",X"10",X"FD",X"86",X"07",X"DD",X"BE",X"07",X"38",X"6E",X"18",X"14",
		X"FD",X"7E",X"08",X"B7",X"20",X"0E",X"78",X"DD",X"86",X"0E",X"C6",X"10",X"DD",X"86",X"07",X"FD",
		X"BE",X"07",X"38",X"58",X"DD",X"7E",X"03",X"FD",X"BE",X"03",X"38",X"50",X"FD",X"7E",X"03",X"BA",
		X"30",X"4A",X"57",X"DD",X"E5",X"DD",X"21",X"66",X"F2",X"DD",X"36",X"00",X"10",X"FD",X"7E",X"05",
		X"D6",X"04",X"DD",X"77",X"01",X"C6",X"18",X"DD",X"77",X"02",X"DD",X"36",X"03",X"F0",X"DD",X"36",
		X"04",X"00",X"FD",X"22",X"3A",X"F0",X"DD",X"E5",X"DD",X"21",X"5B",X"F2",X"FD",X"21",X"71",X"F2",
		X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"B7",X"20",X"F3",X"DD",X"E1",X"FD",
		X"21",X"71",X"F2",X"CD",X"DE",X"44",X"FD",X"2A",X"3A",X"F0",X"DD",X"E1",X"01",X"23",X"00",X"FD",
		X"09",X"1C",X"C3",X"3D",X"15",X"DD",X"7E",X"05",X"DD",X"86",X"04",X"47",X"7A",X"FE",X"FF",X"28",
		X"5C",X"FD",X"21",X"5B",X"F2",X"CD",X"62",X"45",X"38",X"53",X"FD",X"2A",X"3A",X"F0",X"DD",X"7E",
		X"03",X"3D",X"FD",X"BE",X"03",X"38",X"07",X"DD",X"77",X"03",X"DD",X"36",X"0D",X"04",X"DD",X"36",
		X"0C",X"04",X"FD",X"46",X"04",X"79",X"B7",X"3E",X"01",X"28",X"08",X"ED",X"44",X"CB",X"78",X"20",
		X"06",X"18",X"06",X"CB",X"78",X"20",X"02",X"CB",X"27",X"47",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",
		X"06",X"38",X"16",X"3A",X"01",X"F0",X"C6",X"18",X"DD",X"BE",X"07",X"38",X"0C",X"3A",X"01",X"F0",
		X"D6",X"18",X"DD",X"BE",X"07",X"30",X"02",X"06",X"00",X"78",X"C3",X"EE",X"1A",X"3A",X"15",X"F0",
		X"B7",X"28",X"5A",X"DD",X"7E",X"07",X"C6",X"D0",X"30",X"53",X"FD",X"21",X"5B",X"F2",X"4F",X"06",
		X"00",X"CD",X"B5",X"41",X"DD",X"46",X"05",X"CD",X"62",X"45",X"38",X"3A",X"DD",X"7E",X"0D",X"FE",
		X"04",X"30",X"04",X"DD",X"36",X"0D",X"04",X"DD",X"7E",X"0B",X"D6",X"02",X"DD",X"BE",X"03",X"30",
		X"03",X"DD",X"77",X"03",X"DD",X"36",X"0C",X"04",X"DD",X"7E",X"10",X"CB",X"7F",X"28",X"02",X"ED",
		X"44",X"D6",X"02",X"38",X"03",X"B7",X"20",X"02",X"3E",X"01",X"57",X"79",X"B7",X"7A",X"CA",X"EE",
		X"1A",X"ED",X"44",X"C3",X"EE",X"1A",X"DD",X"7E",X"05",X"DD",X"86",X"04",X"47",X"DD",X"70",X"05",
		X"78",X"DD",X"35",X"0C",X"C2",X"1B",X"1B",X"DD",X"36",X"0C",X"01",X"0E",X"00",X"3A",X"15",X"F0",
		X"B7",X"DD",X"7E",X"02",X"CA",X"8B",X"17",X"E6",X"0F",X"FE",X"05",X"CA",X"29",X"19",X"57",X"3A",
		X"06",X"F0",X"FE",X"02",X"CA",X"29",X"19",X"DD",X"BE",X"09",X"C2",X"29",X"19",X"3A",X"03",X"F0",
		X"E6",X"33",X"C2",X"29",X"19",X"7A",X"FE",X"01",X"DA",X"3E",X"17",X"C2",X"29",X"19",X"3A",X"01",
		X"F0",X"D6",X"34",X"DD",X"BE",X"07",X"DA",X"D0",X"18",X"CD",X"B9",X"1B",X"3A",X"00",X"F0",X"DD",
		X"96",X"05",X"30",X"02",X"ED",X"44",X"FE",X"03",X"DC",X"E2",X"40",X"C3",X"29",X"19",X"DD",X"7E",
		X"1C",X"B7",X"28",X"06",X"DD",X"35",X"1C",X"C3",X"D0",X"18",X"3A",X"01",X"F0",X"DD",X"96",X"07",
		X"30",X"02",X"ED",X"44",X"FE",X"40",X"DA",X"D0",X"18",X"CD",X"B9",X"1B",X"1E",X"00",X"21",X"00",
		X"F0",X"DD",X"7E",X"04",X"CB",X"27",X"CB",X"27",X"DD",X"86",X"05",X"D6",X"08",X"57",X"96",X"30",
		X"02",X"ED",X"44",X"FE",X"05",X"38",X"0E",X"7A",X"C6",X"0C",X"96",X"30",X"02",X"ED",X"44",X"FE",
		X"05",X"D2",X"29",X"19",X"1C",X"CD",X"12",X"41",X"C3",X"29",X"19",X"E6",X"0F",X"FE",X"06",X"38",
		X"57",X"3A",X"03",X"F0",X"E6",X"03",X"20",X"50",X"3A",X"06",X"F0",X"FE",X"02",X"28",X"49",X"DD",
		X"BE",X"09",X"20",X"44",X"21",X"58",X"F0",X"7E",X"B7",X"20",X"17",X"3A",X"01",X"F0",X"D6",X"34",
		X"DD",X"BE",X"07",X"DA",X"D0",X"18",X"3A",X"A0",X"F0",X"FE",X"01",X"CA",X"D0",X"18",X"36",X"01",
		X"18",X"0B",X"FE",X"04",X"38",X"07",X"CA",X"29",X"19",X"0C",X"C3",X"29",X"19",X"3A",X"00",X"F0",
		X"DD",X"BE",X"05",X"CA",X"29",X"19",X"30",X"08",X"0D",X"DD",X"36",X"11",X"20",X"C3",X"29",X"19",
		X"0C",X"DD",X"36",X"11",X"E0",X"C3",X"29",X"19",X"3A",X"55",X"F0",X"57",X"E6",X"60",X"28",X"1E",
		X"CB",X"6A",X"28",X"0D",X"0C",X"DD",X"7E",X"03",X"FE",X"09",X"DA",X"29",X"19",X"0C",X"C3",X"29",
		X"19",X"0D",X"DD",X"7E",X"03",X"FE",X"09",X"DA",X"29",X"19",X"0D",X"C3",X"29",X"19",X"7A",X"CB",
		X"5F",X"20",X"10",X"E6",X"0F",X"FE",X"06",X"38",X"0A",X"3E",X"01",X"20",X"02",X"ED",X"44",X"4F",
		X"C3",X"29",X"19",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"02",X"D2",X"29",X"19",X"57",X"3A",X"06",
		X"F0",X"FE",X"02",X"CA",X"29",X"19",X"DD",X"BE",X"09",X"C2",X"29",X"19",X"3A",X"03",X"F0",X"E6",
		X"13",X"C2",X"29",X"19",X"7A",X"B7",X"CA",X"D0",X"18",X"3A",X"01",X"F0",X"DD",X"96",X"07",X"30",
		X"02",X"ED",X"44",X"FE",X"0A",X"30",X"2F",X"3A",X"00",X"F0",X"DD",X"96",X"05",X"57",X"30",X"02",
		X"ED",X"44",X"FE",X"30",X"30",X"24",X"3A",X"14",X"F0",X"B7",X"3E",X"05",X"28",X"02",X"3E",X"03",
		X"CB",X"7A",X"28",X"02",X"ED",X"44",X"4F",X"DD",X"36",X"0C",X"06",X"DD",X"7E",X"01",X"F6",X"04",
		X"DD",X"77",X"01",X"C3",X"29",X"19",X"FE",X"30",X"30",X"46",X"CD",X"56",X"40",X"DD",X"7E",X"0D",
		X"FE",X"02",X"30",X"3C",X"21",X"82",X"F0",X"56",X"3A",X"01",X"F0",X"DD",X"96",X"07",X"3E",X"00",
		X"28",X"05",X"3C",X"38",X"02",X"ED",X"44",X"82",X"CB",X"7F",X"28",X"02",X"ED",X"44",X"57",X"DD",
		X"7E",X"03",X"BA",X"28",X"13",X"38",X"03",X"3D",X"18",X"0B",X"3C",X"DD",X"BE",X"0B",X"28",X"05",
		X"38",X"03",X"DD",X"7E",X"0B",X"DD",X"77",X"03",X"3A",X"41",X"F0",X"C6",X"02",X"DD",X"77",X"0D",
		X"3A",X"00",X"F0",X"DD",X"86",X"11",X"DD",X"96",X"05",X"28",X"4E",X"F5",X"3A",X"01",X"F0",X"C6",
		X"1C",X"DD",X"BE",X"07",X"30",X"14",X"DD",X"7E",X"10",X"CB",X"7F",X"28",X"0D",X"3A",X"82",X"F0",
		X"B7",X"28",X"07",X"DD",X"77",X"03",X"DD",X"36",X"0D",X"01",X"F1",X"38",X"03",X"0C",X"18",X"03",
		X"0D",X"ED",X"44",X"FE",X"40",X"38",X"0A",X"DD",X"7E",X"11",X"ED",X"44",X"DD",X"77",X"11",X"18",
		X"18",X"FE",X"04",X"38",X"14",X"DD",X"7E",X"06",X"FE",X"27",X"20",X"0D",X"3A",X"01",X"F0",X"DD",
		X"96",X"0E",X"DD",X"BE",X"07",X"38",X"02",X"CB",X"21",X"DD",X"71",X"04",X"78",X"C3",X"1B",X"1B",
		X"E6",X"04",X"28",X"6F",X"78",X"E6",X"02",X"20",X"5E",X"DD",X"7E",X"0C",X"FE",X"80",X"30",X"08",
		X"3D",X"DD",X"77",X"0C",X"28",X"51",X"18",X"5B",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"05",X"30",
		X"52",X"DD",X"35",X"22",X"20",X"4D",X"DD",X"36",X"22",X"06",X"DD",X"7E",X"21",X"3C",X"E6",X"03",
		X"DD",X"77",X"21",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"01",X"20",X"03",X"DD",X"86",X"16",X"21",
		X"04",X"1C",X"CB",X"27",X"85",X"30",X"01",X"24",X"6F",X"5E",X"23",X"56",X"D5",X"E1",X"DD",X"7E",
		X"21",X"CB",X"27",X"85",X"30",X"01",X"24",X"6F",X"7E",X"DD",X"77",X"06",X"3C",X"DD",X"77",X"1D",
		X"23",X"7E",X"DD",X"77",X"1E",X"18",X"0C",X"DD",X"36",X"0C",X"01",X"DD",X"7E",X"01",X"EE",X"04",
		X"DD",X"77",X"01",X"78",X"E6",X"08",X"CA",X"0F",X"1B",X"DD",X"7E",X"16",X"47",X"B7",X"20",X"74",
		X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"05",X"38",X"20",X"FD",X"21",X"68",X"F8",X"FD",X"36",X"00",
		X"00",X"DD",X"36",X"16",X"7F",X"DD",X"7E",X"18",X"B7",X"CA",X"90",X"1A",X"67",X"DD",X"6E",X"17",
		X"36",X"00",X"DD",X"36",X"18",X"00",X"C3",X"90",X"1A",X"FE",X"02",X"20",X"09",X"DD",X"36",X"18",
		X"00",X"3E",X"80",X"47",X"18",X"45",X"DD",X"7E",X"18",X"B7",X"28",X"06",X"67",X"DD",X"6E",X"17",
		X"18",X"0F",X"CD",X"EF",X"1B",X"DA",X"90",X"1A",X"FD",X"E5",X"E1",X"DD",X"75",X"17",X"DD",X"74",
		X"18",X"0E",X"17",X"CD",X"4E",X"3D",X"DD",X"7E",X"02",X"E6",X"0F",X"CB",X"27",X"21",X"DD",X"1B",
		X"85",X"30",X"01",X"24",X"6F",X"7E",X"DD",X"77",X"19",X"23",X"7E",X"DD",X"77",X"1A",X"DD",X"36",
		X"1B",X"38",X"18",X"5D",X"FE",X"7F",X"38",X"23",X"CA",X"90",X"1A",X"E6",X"70",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"21",X"E7",X"1B",X"85",X"30",X"01",X"24",X"6F",X"7E",X"DD",X"77",
		X"06",X"78",X"C6",X"02",X"F6",X"80",X"DD",X"77",X"16",X"18",X"45",X"DD",X"35",X"1C",X"20",X"40",
		X"FE",X"04",X"20",X"11",X"DD",X"35",X"19",X"DD",X"36",X"1B",X"4B",X"DD",X"7E",X"1A",X"C6",X"03",
		X"DD",X"77",X"1A",X"18",X"1C",X"FE",X"08",X"20",X"0B",X"DD",X"36",X"1B",X"4B",X"0E",X"18",X"CD",
		X"4E",X"3D",X"18",X"0D",X"FE",X"0C",X"20",X"06",X"DD",X"36",X"1B",X"4B",X"18",X"03",X"DD",X"34",
		X"1B",X"DD",X"36",X"1C",X"04",X"78",X"3C",X"FE",X"10",X"38",X"02",X"3E",X"0C",X"DD",X"77",X"16",
		X"DD",X"7E",X"1F",X"B7",X"20",X"11",X"DD",X"35",X"20",X"20",X"0C",X"DD",X"7E",X"01",X"F6",X"03",
		X"DD",X"77",X"01",X"DD",X"36",X"1F",X"10",X"DD",X"35",X"0C",X"20",X"63",X"3A",X"82",X"F0",X"FE",
		X"04",X"DD",X"7E",X"03",X"38",X"09",X"21",X"40",X"F0",X"86",X"CB",X"3F",X"DD",X"77",X"03",X"B7",
		X"28",X"2C",X"CD",X"E7",X"3C",X"47",X"E6",X"07",X"3C",X"DD",X"77",X"0C",X"DD",X"7E",X"03",X"0E",
		X"03",X"FE",X"04",X"30",X"02",X"CB",X"39",X"78",X"A1",X"CB",X"58",X"28",X"02",X"ED",X"44",X"FE",
		X"02",X"38",X"0B",X"3A",X"15",X"F0",X"B7",X"20",X"05",X"0E",X"26",X"CD",X"4E",X"3D",X"47",X"DD",
		X"7E",X"04",X"CB",X"7F",X"20",X"0C",X"CB",X"78",X"20",X"05",X"B8",X"28",X"0F",X"38",X"0C",X"3D",
		X"18",X"0A",X"CB",X"78",X"28",X"05",X"B8",X"28",X"03",X"30",X"F4",X"3C",X"DD",X"77",X"04",X"DD",
		X"7E",X"03",X"B7",X"DD",X"7E",X"05",X"28",X"03",X"DD",X"86",X"04",X"FE",X"06",X"38",X"0A",X"FE",
		X"FA",X"30",X"06",X"DD",X"77",X"05",X"C3",X"B7",X"1B",X"CD",X"32",X"3F",X"DD",X"7E",X"02",X"E6",
		X"0F",X"20",X"21",X"3A",X"06",X"F0",X"DD",X"BE",X"09",X"C2",X"B7",X"1B",X"21",X"59",X"B9",X"CD",
		X"EE",X"3D",X"3A",X"8E",X"F3",X"FE",X"02",X"38",X"63",X"21",X"E7",X"F0",X"7E",X"B7",X"20",X"5C",
		X"36",X"80",X"18",X"58",X"FE",X"06",X"38",X"42",X"3A",X"06",X"F0",X"DD",X"BE",X"09",X"20",X"57",
		X"3A",X"0A",X"F0",X"B7",X"20",X"51",X"3A",X"03",X"F0",X"B7",X"20",X"46",X"3A",X"06",X"F0",X"FE",
		X"02",X"30",X"3F",X"21",X"28",X"F0",X"3A",X"8E",X"F3",X"3C",X"CB",X"27",X"C6",X"08",X"86",X"77",
		X"3A",X"5E",X"F0",X"B7",X"28",X"2C",X"AF",X"32",X"5E",X"F0",X"3A",X"5D",X"F0",X"B7",X"20",X"22",
		X"3A",X"12",X"F0",X"EE",X"04",X"32",X"12",X"F0",X"18",X"18",X"FE",X"01",X"20",X"BA",X"3A",X"06",
		X"F0",X"DD",X"BE",X"09",X"20",X"11",X"21",X"52",X"B9",X"CD",X"EE",X"3D",X"3A",X"0A",X"F0",X"B7",
		X"20",X"05",X"0E",X"17",X"CD",X"4E",X"3D",X"D1",X"C9",X"3A",X"00",X"F0",X"DD",X"86",X"11",X"DD",
		X"96",X"05",X"20",X"0A",X"DD",X"7E",X"11",X"ED",X"44",X"DD",X"77",X"11",X"18",X"EB",X"0E",X"02",
		X"30",X"04",X"0E",X"FE",X"ED",X"44",X"FE",X"04",X"30",X"02",X"CB",X"29",X"C9",X"01",X"13",X"02",
		X"0A",X"00",X"00",X"02",X"06",X"02",X"0A",X"4F",X"24",X"50",X"24",X"4F",X"24",X"50",X"24",X"0E",
		X"06",X"FD",X"21",X"DC",X"F8",X"11",X"04",X"00",X"FD",X"7E",X"00",X"B7",X"C8",X"FD",X"19",X"0D",
		X"20",X"F6",X"37",X"C9",X"10",X"1C",X"18",X"1C",X"20",X"1C",X"30",X"1C",X"38",X"1C",X"28",X"1C",
		X"25",X"00",X"C9",X"FE",X"25",X"00",X"DE",X"02",X"7C",X"00",X"CB",X"00",X"7C",X"00",X"CD",X"00",
		X"24",X"00",X"4F",X"00",X"24",X"00",X"50",X"00",X"27",X"00",X"CF",X"00",X"27",X"00",X"D1",X"00",
		X"23",X"00",X"DC",X"00",X"23",X"00",X"DD",X"00",X"2C",X"00",X"E0",X"00",X"2C",X"00",X"E2",X"00",
		X"3A",X"03",X"F0",X"57",X"E6",X"10",X"C0",X"7A",X"E6",X"01",X"C2",X"D3",X"66",X"7A",X"E6",X"02",
		X"28",X"37",X"21",X"05",X"F0",X"35",X"20",X"14",X"36",X"04",X"21",X"02",X"F0",X"3A",X"A1",X"F0",
		X"CB",X"7F",X"28",X"03",X"34",X"18",X"01",X"35",X"7E",X"E6",X"07",X"77",X"3A",X"01",X"F0",X"FE",
		X"30",X"38",X"01",X"3D",X"3D",X"32",X"01",X"F0",X"21",X"00",X"F0",X"3A",X"A1",X"F0",X"B7",X"20",
		X"05",X"3E",X"02",X"32",X"A1",X"F0",X"86",X"77",X"C9",X"7A",X"E6",X"04",X"28",X"18",X"0E",X"26",
		X"CD",X"4E",X"3D",X"21",X"27",X"F0",X"35",X"20",X"0D",X"3A",X"03",X"F0",X"EE",X"04",X"32",X"03",
		X"F0",X"21",X"02",X"F0",X"36",X"08",X"2A",X"81",X"F0",X"E5",X"C1",X"29",X"29",X"09",X"3A",X"15",
		X"F0",X"B7",X"28",X"02",X"09",X"09",X"3E",X"D0",X"94",X"32",X"01",X"F0",X"FE",X"D0",X"C8",X"3A",
		X"0A",X"F0",X"B7",X"C0",X"3A",X"82",X"F0",X"B7",X"C8",X"47",X"ED",X"44",X"4F",X"3A",X"15",X"F0",
		X"57",X"21",X"19",X"F0",X"1E",X"00",X"3A",X"18",X"F0",X"B6",X"28",X"07",X"1C",X"7E",X"B7",X"20",
		X"02",X"1C",X"1C",X"3A",X"A1",X"F0",X"ED",X"44",X"CB",X"42",X"28",X"02",X"CB",X"2F",X"21",X"00",
		X"F0",X"CB",X"7F",X"28",X"0B",X"B9",X"30",X"01",X"79",X"86",X"38",X"0B",X"3E",X"10",X"18",X"65",
		X"B8",X"38",X"01",X"78",X"86",X"38",X"5C",X"CB",X"43",X"28",X"0E",X"CB",X"4B",X"16",X"2A",X"20",
		X"02",X"16",X"BA",X"BA",X"30",X"1F",X"7A",X"18",X"4C",X"FE",X"10",X"30",X"18",X"3A",X"03",X"F0",
		X"E6",X"04",X"28",X"D8",X"F6",X"02",X"32",X"03",X"F0",X"3A",X"A1",X"F0",X"ED",X"44",X"32",X"A1",
		X"F0",X"CD",X"AF",X"7D",X"C9",X"CB",X"43",X"28",X"0E",X"CB",X"4B",X"16",X"3A",X"20",X"02",X"16",
		X"C6",X"BA",X"38",X"21",X"7A",X"18",X"1E",X"FE",X"F0",X"38",X"1A",X"3A",X"03",X"F0",X"E6",X"04",
		X"28",X"11",X"F6",X"02",X"32",X"03",X"F0",X"3A",X"A1",X"F0",X"ED",X"44",X"32",X"A1",X"F0",X"CD",
		X"AF",X"7D",X"C9",X"3E",X"F0",X"77",X"3A",X"03",X"F0",X"E6",X"40",X"C0",X"7B",X"B7",X"C0",X"21",
		X"02",X"F0",X"3A",X"A1",X"F0",X"06",X"07",X"CB",X"7F",X"28",X"04",X"06",X"00",X"ED",X"44",X"FE",
		X"07",X"30",X"03",X"36",X"08",X"C9",X"70",X"0E",X"26",X"CB",X"42",X"CC",X"4E",X"3D",X"C9",X"AF",
		X"32",X"09",X"F0",X"32",X"56",X"F0",X"5F",X"21",X"01",X"F0",X"4E",X"06",X"00",X"CD",X"5A",X"4B",
		X"3A",X"00",X"F0",X"C6",X"04",X"47",X"DD",X"7E",X"00",X"57",X"21",X"56",X"F0",X"B6",X"77",X"7A",
		X"E6",X"0F",X"57",X"FE",X"06",X"28",X"09",X"FE",X"0E",X"28",X"05",X"DD",X"7E",X"01",X"B8",X"D0",
		X"7A",X"CB",X"27",X"82",X"21",X"D1",X"1D",X"85",X"30",X"01",X"24",X"6F",X"78",X"DD",X"96",X"01",
		X"E9",X"C3",X"01",X"1E",X"C3",X"0F",X"1E",X"C3",X"26",X"1E",X"C3",X"36",X"1E",X"C3",X"5F",X"1E",
		X"C3",X"C7",X"1E",X"C3",X"F1",X"1E",X"C3",X"0B",X"1F",X"C3",X"34",X"1F",X"C3",X"59",X"1F",X"C3",
		X"7E",X"1F",X"C3",X"34",X"1F",X"C3",X"59",X"1F",X"C3",X"7E",X"1F",X"C3",X"AF",X"1F",X"C3",X"E9",
		X"1F",X"F5",X"3A",X"15",X"F0",X"B7",X"20",X"03",X"F1",X"18",X"2B",X"F1",X"C3",X"7E",X"1F",X"D6",
		X"14",X"38",X"6C",X"C6",X"10",X"DD",X"96",X"02",X"DA",X"A1",X"1E",X"DD",X"96",X"03",X"DA",X"A1",
		X"1E",X"D6",X"14",X"38",X"5A",X"C9",X"D6",X"14",X"38",X"55",X"C6",X"10",X"DD",X"96",X"02",X"38",
		X"70",X"D6",X"14",X"38",X"4A",X"C9",X"D6",X"14",X"38",X"45",X"C6",X"10",X"DD",X"96",X"02",X"38",
		X"60",X"D6",X"12",X"38",X"3A",X"D6",X"10",X"38",X"7C",X"C6",X"02",X"DD",X"96",X"03",X"38",X"75",
		X"D6",X"12",X"38",X"2B",X"C6",X"10",X"D6",X"50",X"38",X"43",X"D6",X"14",X"38",X"21",X"C9",X"D6",
		X"10",X"38",X"1C",X"C6",X"0E",X"DD",X"96",X"02",X"38",X"37",X"D6",X"0E",X"38",X"11",X"DD",X"96",
		X"03",X"38",X"0C",X"C6",X"0E",X"DD",X"96",X"02",X"38",X"23",X"D6",X"14",X"38",X"01",X"C9",X"3A",
		X"15",X"F0",X"B7",X"28",X"11",X"3A",X"82",X"F0",X"FE",X"04",X"38",X"0A",X"3A",X"03",X"F0",X"F6",
		X"40",X"32",X"03",X"F0",X"18",X"0D",X"21",X"09",X"F0",X"36",X"01",X"18",X"06",X"16",X"01",X"18",
		X"02",X"16",X"00",X"7B",X"B7",X"28",X"13",X"3A",X"09",X"F0",X"B7",X"20",X"0B",X"3A",X"03",X"F0",
		X"E6",X"40",X"20",X"04",X"7A",X"32",X"06",X"F0",X"37",X"C9",X"1C",X"3A",X"04",X"F0",X"D6",X"04",
		X"81",X"4F",X"C3",X"9B",X"1D",X"3F",X"C9",X"D6",X"14",X"38",X"B4",X"C6",X"10",X"DD",X"96",X"02",
		X"38",X"CF",X"D6",X"12",X"38",X"A9",X"D6",X"10",X"38",X"EB",X"C6",X"02",X"DD",X"96",X"03",X"38",
		X"E4",X"D6",X"12",X"38",X"9A",X"C6",X"10",X"DD",X"96",X"02",X"38",X"B1",X"D6",X"14",X"38",X"8F",
		X"C9",X"D6",X"20",X"38",X"D0",X"DD",X"96",X"02",X"38",X"CB",X"D6",X"10",X"38",X"81",X"C6",X"0E",
		X"DD",X"96",X"03",X"38",X"98",X"D6",X"10",X"DA",X"7F",X"1E",X"C9",X"D6",X"10",X"DA",X"7F",X"1E",
		X"C6",X"0E",X"DD",X"96",X"02",X"38",X"8A",X"D6",X"10",X"DA",X"7F",X"1E",X"C9",X"78",X"D6",X"82",
		X"38",X"A3",X"D6",X"14",X"DA",X"7F",X"1E",X"C6",X"10",X"D6",X"50",X"DA",X"A1",X"1E",X"D6",X"14",
		X"DA",X"7F",X"1E",X"C9",X"D6",X"10",X"DA",X"7F",X"1E",X"C6",X"0E",X"DD",X"96",X"02",X"DA",X"A1",
		X"1E",X"D6",X"0E",X"DA",X"7F",X"1E",X"D6",X"10",X"DA",X"7F",X"1E",X"C6",X"0E",X"DD",X"96",X"03",
		X"DA",X"9D",X"1E",X"D6",X"14",X"DA",X"7F",X"1E",X"C9",X"D6",X"10",X"DA",X"7F",X"1E",X"C6",X"0E",
		X"DD",X"96",X"02",X"DA",X"A1",X"1E",X"D6",X"0E",X"DA",X"7F",X"1E",X"D6",X"20",X"DA",X"7F",X"1E",
		X"C6",X"0E",X"DD",X"96",X"03",X"DA",X"9D",X"1E",X"D6",X"14",X"DA",X"7F",X"1E",X"C9",X"D6",X"14",
		X"DA",X"7F",X"1E",X"C6",X"10",X"DD",X"96",X"02",X"DA",X"A1",X"1E",X"D6",X"12",X"DA",X"7F",X"1E",
		X"D6",X"10",X"DA",X"C5",X"1E",X"C6",X"02",X"D6",X"20",X"DA",X"C5",X"1E",X"D6",X"12",X"DA",X"7F",
		X"1E",X"C6",X"10",X"DD",X"96",X"03",X"DA",X"9D",X"1E",X"D6",X"14",X"DA",X"7F",X"1E",X"C9",X"DD",
		X"7E",X"01",X"B7",X"C8",X"78",X"D6",X"34",X"D8",X"D6",X"14",X"DA",X"7F",X"1E",X"C6",X"10",X"D6",
		X"30",X"DA",X"A1",X"1E",X"D6",X"12",X"DA",X"7F",X"1E",X"D6",X"10",X"DA",X"C5",X"1E",X"C6",X"02",
		X"DD",X"96",X"01",X"DA",X"C5",X"1E",X"D6",X"12",X"DA",X"7F",X"1E",X"C6",X"10",X"DD",X"96",X"02",
		X"DA",X"9D",X"1E",X"D6",X"14",X"DA",X"9D",X"1E",X"C9",X"3A",X"15",X"F0",X"B7",X"3A",X"00",X"F0",
		X"28",X"1F",X"FE",X"80",X"38",X"14",X"3A",X"03",X"F0",X"E6",X"03",X"20",X"0D",X"3A",X"19",X"F0",
		X"B7",X"20",X"07",X"3C",X"32",X"06",X"F0",X"32",X"19",X"F0",X"78",X"DD",X"96",X"01",X"C3",X"7E",
		X"1F",X"FE",X"60",X"30",X"14",X"3A",X"03",X"F0",X"E6",X"03",X"20",X"0D",X"3A",X"18",X"F0",X"B7",
		X"20",X"07",X"32",X"06",X"F0",X"3C",X"32",X"18",X"F0",X"78",X"DD",X"96",X"01",X"C3",X"36",X"1E",
		X"3A",X"0A",X"F0",X"B7",X"37",X"C0",X"21",X"15",X"F0",X"3A",X"16",X"F0",X"BE",X"37",X"C0",X"D5",
		X"FD",X"E5",X"DD",X"E5",X"1E",X"00",X"DD",X"4E",X"07",X"06",X"00",X"CD",X"5A",X"4B",X"FD",X"E1",
		X"DD",X"7E",X"00",X"32",X"54",X"F0",X"E6",X"0F",X"6F",X"CB",X"27",X"85",X"21",X"68",X"20",X"85",
		X"30",X"01",X"24",X"6F",X"FD",X"7E",X"05",X"E9",X"C3",X"98",X"20",X"C3",X"A3",X"20",X"C3",X"BF",
		X"20",X"C3",X"D5",X"20",X"C3",X"EE",X"20",X"C3",X"34",X"21",X"C3",X"62",X"21",X"C3",X"81",X"21",
		X"C3",X"D5",X"20",X"C3",X"EF",X"21",X"C3",X"39",X"22",X"C3",X"8F",X"22",X"C3",X"BC",X"22",X"C3",
		X"E9",X"22",X"C3",X"20",X"23",X"C3",X"43",X"23",X"F5",X"3A",X"15",X"F0",X"B7",X"C2",X"40",X"22",
		X"F1",X"18",X"32",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"38",X"67",X"C6",X"10",X"DD",
		X"96",X"02",X"38",X"60",X"DD",X"96",X"03",X"38",X"5B",X"D6",X"10",X"38",X"57",X"18",X"6D",X"DD",
		X"96",X"01",X"38",X"67",X"D6",X"10",X"38",X"4C",X"C6",X"10",X"DD",X"96",X"02",X"38",X"45",X"D6",
		X"10",X"38",X"41",X"18",X"57",X"D6",X"82",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C6",
		X"10",X"D6",X"50",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C3",X"2C",X"21",X"DD",X"96",
		X"01",X"38",X"38",X"D6",X"10",X"38",X"1D",X"C6",X"10",X"DD",X"96",X"02",X"38",X"16",X"D6",X"10",
		X"38",X"12",X"DD",X"96",X"03",X"38",X"0D",X"C6",X"10",X"DD",X"96",X"02",X"38",X"06",X"D6",X"10",
		X"38",X"02",X"18",X"18",X"7B",X"B7",X"28",X"03",X"37",X"18",X"11",X"1C",X"06",X"00",X"FD",X"7E",
		X"0E",X"81",X"4F",X"30",X"01",X"04",X"FD",X"E5",X"C3",X"4B",X"20",X"3F",X"FD",X"E5",X"DD",X"E1",
		X"FD",X"E1",X"D1",X"C9",X"DD",X"96",X"01",X"38",X"F2",X"D6",X"10",X"38",X"D7",X"C6",X"10",X"DD",
		X"96",X"02",X"38",X"D0",X"D6",X"10",X"38",X"CC",X"D6",X"10",X"38",X"DF",X"DD",X"96",X"03",X"38",
		X"DA",X"D6",X"10",X"38",X"BF",X"C6",X"10",X"DD",X"96",X"02",X"38",X"B8",X"D6",X"10",X"38",X"B4",
		X"18",X"CA",X"C6",X"10",X"DD",X"96",X"01",X"38",X"AB",X"D6",X"20",X"38",X"A7",X"DD",X"96",X"02",
		X"38",X"B9",X"D6",X"10",X"38",X"9E",X"DD",X"96",X"03",X"38",X"99",X"D6",X"10",X"38",X"95",X"18",
		X"AB",X"DD",X"96",X"01",X"38",X"A5",X"D6",X"10",X"38",X"8A",X"C6",X"10",X"DD",X"96",X"02",X"38",
		X"83",X"D6",X"10",X"DA",X"14",X"21",X"DD",X"96",X"03",X"38",X"90",X"C3",X"14",X"21",X"F5",X"3A",
		X"15",X"F0",X"B7",X"28",X"21",X"F1",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"14",
		X"21",X"C6",X"10",X"DD",X"96",X"02",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"D6",X"10",
		X"DA",X"14",X"21",X"C3",X"2C",X"21",X"F1",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"DA",
		X"2B",X"21",X"C6",X"10",X"DD",X"96",X"02",X"DA",X"2B",X"21",X"D6",X"20",X"DA",X"14",X"21",X"C6",
		X"10",X"DD",X"96",X"03",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C3",X"2C",X"21",X"F5",
		X"3A",X"15",X"F0",X"B7",X"28",X"1C",X"F1",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"DA",
		X"14",X"21",X"C6",X"10",X"DD",X"96",X"02",X"DA",X"14",X"21",X"D6",X"30",X"DA",X"14",X"21",X"C3",
		X"2C",X"21",X"F1",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"2B",X"21",X"C6",X"10",
		X"DD",X"96",X"02",X"DA",X"2B",X"21",X"D6",X"30",X"DA",X"14",X"21",X"DD",X"96",X"03",X"DA",X"14",
		X"21",X"D6",X"10",X"DA",X"14",X"21",X"C3",X"2C",X"21",X"F5",X"3A",X"15",X"F0",X"B7",X"28",X"21",
		X"F1",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C6",X"10",X"DD",X"96",
		X"02",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"D6",X"30",X"DA",X"2B",X"21",X"C3",X"2C",
		X"21",X"F1",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"2B",X"21",X"C6",X"10",X"DD",
		X"96",X"02",X"DA",X"2B",X"21",X"D6",X"30",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C6",
		X"10",X"DD",X"96",X"03",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C3",X"2C",X"21",X"DD",
		X"96",X"01",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C6",X"10",X"DD",X"96",X"02",X"DA",
		X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C6",X"10",X"DD",X"96",
		X"03",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C3",X"2C",X"21",X"DD",X"96",X"01",X"DA",
		X"2B",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C6",X"10",X"DD",X"96",X"02",X"DA",X"14",X"21",X"D6",
		X"10",X"DA",X"14",X"21",X"D6",X"20",X"DA",X"14",X"21",X"C6",X"10",X"DD",X"96",X"03",X"DA",X"14",
		X"21",X"D6",X"10",X"DA",X"14",X"21",X"C3",X"2C",X"21",X"DD",X"96",X"01",X"DA",X"2B",X"21",X"D6",
		X"10",X"DA",X"14",X"21",X"C6",X"10",X"DD",X"96",X"02",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",
		X"21",X"D6",X"10",X"DA",X"2B",X"21",X"D6",X"20",X"DA",X"2B",X"21",X"D6",X"10",X"DA",X"14",X"21",
		X"C6",X"10",X"DD",X"96",X"03",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",X"C3",X"2C",X"21",
		X"DD",X"7E",X"01",X"B7",X"CA",X"2C",X"21",X"FD",X"7E",X"05",X"D6",X"34",X"DA",X"2B",X"21",X"D6",
		X"10",X"DA",X"14",X"21",X"C6",X"10",X"D6",X"30",X"DA",X"14",X"21",X"D6",X"10",X"DA",X"14",X"21",
		X"C3",X"2C",X"21",X"F5",X"3A",X"15",X"F0",X"B7",X"C2",X"40",X"22",X"F1",X"C3",X"D5",X"20",X"3A",
		X"25",X"F0",X"B7",X"C0",X"16",X"00",X"DD",X"21",X"78",X"F8",X"21",X"3B",X"F1",X"01",X"04",X"00",
		X"DD",X"7E",X"00",X"B7",X"28",X"20",X"CD",X"AB",X"45",X"38",X"17",X"7E",X"B7",X"28",X"13",X"35",
		X"DD",X"7E",X"03",X"D6",X"10",X"DD",X"77",X"03",X"DD",X"7E",X"01",X"EE",X"20",X"DD",X"77",X"01",
		X"18",X"09",X"DD",X"36",X"00",X"00",X"DD",X"E5",X"FD",X"E1",X"5A",X"DD",X"09",X"23",X"14",X"7A",
		X"FE",X"06",X"20",X"CC",X"DD",X"21",X"74",X"F8",X"DD",X"7E",X"00",X"B7",X"28",X"28",X"DD",X"7E",
		X"01",X"EE",X"20",X"DD",X"77",X"01",X"FD",X"77",X"01",X"FD",X"36",X"02",X"0F",X"DD",X"7E",X"00",
		X"FD",X"77",X"00",X"DD",X"7E",X"03",X"D6",X"10",X"FD",X"77",X"03",X"21",X"3B",X"F1",X"7B",X"85",
		X"30",X"01",X"24",X"6F",X"36",X"05",X"3A",X"11",X"F0",X"B7",X"20",X"16",X"DB",X"01",X"2F",X"E6",
		X"10",X"B7",X"28",X"2E",X"3A",X"03",X"F0",X"E6",X"13",X"20",X"27",X"3A",X"12",X"F0",X"E6",X"01",
		X"28",X"20",X"3A",X"10",X"F0",X"FE",X"03",X"28",X"0A",X"3E",X"03",X"32",X"10",X"F0",X"0E",X"22",
		X"CD",X"4E",X"3D",X"3A",X"00",X"F0",X"DD",X"77",X"00",X"3A",X"01",X"F0",X"D6",X"10",X"DD",X"77",
		X"03",X"C9",X"3A",X"10",X"F0",X"B7",X"C8",X"3D",X"32",X"10",X"F0",X"AF",X"DD",X"77",X"00",X"0E",
		X"23",X"CD",X"4E",X"3D",X"C9",X"3A",X"03",X"F0",X"E6",X"80",X"C0",X"3A",X"58",X"F0",X"FE",X"01",
		X"38",X"32",X"3D",X"47",X"CB",X"27",X"80",X"21",X"A2",X"24",X"85",X"30",X"01",X"24",X"6F",X"E5",
		X"CD",X"35",X"24",X"E1",X"E9",X"DD",X"2A",X"5F",X"F0",X"DD",X"7E",X"01",X"E6",X"03",X"C0",X"21",
		X"59",X"F0",X"35",X"C0",X"36",X"06",X"DD",X"7E",X"06",X"06",X"D3",X"B8",X"20",X"02",X"06",X"29",
		X"DD",X"70",X"06",X"C9",X"3A",X"57",X"F0",X"B7",X"20",X"2B",X"3A",X"60",X"F0",X"B7",X"28",X"05",
		X"CD",X"35",X"24",X"18",X"20",X"DB",X"01",X"2F",X"E6",X"04",X"C8",X"3A",X"57",X"F0",X"B7",X"C0",
		X"3A",X"5E",X"F0",X"B7",X"C8",X"3E",X"01",X"32",X"57",X"F0",X"32",X"5D",X"F0",X"AF",X"32",X"5C",
		X"F0",X"32",X"5E",X"F0",X"C9",X"21",X"5D",X"F0",X"35",X"C0",X"36",X"10",X"3A",X"5C",X"F0",X"EE",
		X"04",X"32",X"5C",X"F0",X"C9",X"AF",X"32",X"5C",X"F0",X"32",X"58",X"F0",X"3E",X"29",X"DD",X"77",
		X"06",X"C9",X"C3",X"C0",X"24",X"C3",X"F8",X"24",X"C3",X"9F",X"25",X"C3",X"F6",X"25",X"C3",X"16",
		X"26",X"C3",X"87",X"26",X"C3",X"CD",X"26",X"C3",X"E3",X"26",X"C3",X"04",X"27",X"C3",X"44",X"27",
		X"DD",X"7E",X"01",X"E6",X"0A",X"20",X"CE",X"3A",X"A0",X"F0",X"FE",X"01",X"28",X"C7",X"FD",X"21",
		X"68",X"F8",X"DD",X"7E",X"05",X"FD",X"77",X"00",X"FD",X"36",X"02",X"2B",X"DD",X"7E",X"07",X"C6",
		X"1C",X"FD",X"77",X"03",X"DD",X"36",X"0B",X"0A",X"21",X"58",X"F0",X"36",X"02",X"DD",X"7E",X"01",
		X"E6",X"FE",X"DD",X"77",X"01",X"C3",X"85",X"24",X"DD",X"7E",X"01",X"E6",X"0A",X"20",X"96",X"FD",
		X"21",X"68",X"F8",X"3A",X"03",X"F0",X"E6",X"03",X"20",X"2C",X"3A",X"A0",X"F0",X"FE",X"01",X"28",
		X"25",X"DD",X"7E",X"08",X"FE",X"01",X"38",X"17",X"28",X"1C",X"DD",X"7E",X"07",X"FE",X"E2",X"38",
		X"15",X"C6",X"20",X"FD",X"77",X"03",X"DD",X"7E",X"05",X"FD",X"77",X"00",X"C3",X"85",X"24",X"DD",
		X"7E",X"07",X"FE",X"D7",X"38",X"0A",X"AF",X"FD",X"77",X"00",X"32",X"58",X"F0",X"C3",X"85",X"24",
		X"C6",X"20",X"FD",X"77",X"03",X"DD",X"7E",X"05",X"FD",X"77",X"00",X"47",X"3A",X"00",X"F0",X"90",
		X"CB",X"7F",X"28",X"02",X"ED",X"44",X"FE",X"03",X"30",X"32",X"DD",X"7E",X"07",X"C6",X"18",X"21",
		X"01",X"F0",X"96",X"30",X"02",X"ED",X"44",X"FE",X"08",X"D2",X"85",X"24",X"3E",X"10",X"32",X"03",
		X"F0",X"21",X"7A",X"F3",X"7E",X"32",X"7B",X"F3",X"36",X"00",X"21",X"81",X"F0",X"36",X"00",X"21",
		X"58",X"F0",X"36",X"03",X"21",X"5A",X"F0",X"36",X"20",X"C3",X"85",X"24",X"FE",X"10",X"DA",X"85",
		X"24",X"DD",X"7E",X"07",X"C6",X"20",X"21",X"01",X"F0",X"96",X"30",X"9A",X"C3",X"85",X"24",X"FD",
		X"21",X"68",X"F8",X"DD",X"7E",X"03",X"FE",X"0C",X"38",X"04",X"3D",X"DD",X"77",X"03",X"32",X"82",
		X"F0",X"DD",X"7E",X"09",X"32",X"06",X"F0",X"3A",X"5A",X"F0",X"D6",X"04",X"FE",X"08",X"28",X"18",
		X"32",X"5A",X"F0",X"DD",X"86",X"07",X"FD",X"77",X"03",X"32",X"01",X"F0",X"DD",X"7E",X"05",X"FD",
		X"77",X"00",X"32",X"00",X"F0",X"C3",X"85",X"24",X"AF",X"FD",X"77",X"00",X"32",X"00",X"F0",X"3E",
		X"10",X"32",X"03",X"F0",X"21",X"5A",X"F0",X"36",X"08",X"21",X"58",X"F0",X"36",X"04",X"21",X"A6",
		X"F0",X"36",X"11",X"C3",X"85",X"24",X"DD",X"7E",X"03",X"32",X"82",X"F0",X"DD",X"7E",X"09",X"32",
		X"06",X"F0",X"21",X"09",X"F4",X"36",X"02",X"21",X"5A",X"F0",X"35",X"C2",X"85",X"24",X"21",X"58",
		X"F0",X"36",X"05",X"C3",X"85",X"24",X"DD",X"7E",X"01",X"E6",X"02",X"20",X"1E",X"DD",X"7E",X"05",
		X"FE",X"F0",X"30",X"17",X"DD",X"7E",X"03",X"B7",X"20",X"05",X"3E",X"02",X"DD",X"77",X"03",X"32",
		X"82",X"F0",X"DD",X"7E",X"09",X"32",X"06",X"F0",X"C3",X"85",X"24",X"AF",X"DD",X"77",X"04",X"DD",
		X"77",X"03",X"32",X"82",X"F0",X"06",X"00",X"0E",X"D0",X"FD",X"21",X"5B",X"F2",X"CD",X"B5",X"41",
		X"DD",X"7E",X"09",X"B7",X"28",X"0B",X"FD",X"7E",X"02",X"B7",X"28",X"05",X"FD",X"7E",X"03",X"18",
		X"0A",X"FD",X"7E",X"01",X"FE",X"60",X"30",X"03",X"FD",X"7E",X"03",X"C6",X"03",X"32",X"07",X"F0",
		X"DD",X"BE",X"05",X"3E",X"00",X"28",X"05",X"3C",X"30",X"02",X"ED",X"44",X"32",X"5A",X"F0",X"21",
		X"58",X"F0",X"36",X"06",X"C3",X"85",X"24",X"DD",X"7E",X"07",X"C6",X"02",X"DD",X"77",X"07",X"FE",
		X"A0",X"30",X"17",X"3A",X"5A",X"F0",X"DD",X"86",X"05",X"DD",X"77",X"05",X"21",X"07",X"F0",X"BE",
		X"C2",X"85",X"24",X"AF",X"32",X"5A",X"F0",X"C3",X"85",X"24",X"DD",X"7E",X"05",X"32",X"00",X"F0",
		X"21",X"01",X"F0",X"36",X"AC",X"FD",X"21",X"68",X"F8",X"FD",X"77",X"00",X"FD",X"36",X"03",X"B0",
		X"21",X"58",X"F0",X"36",X"07",X"21",X"5A",X"F0",X"36",X"10",X"C3",X"85",X"24",X"FD",X"21",X"68",
		X"F8",X"FD",X"34",X"03",X"21",X"5A",X"F0",X"35",X"C2",X"85",X"24",X"21",X"58",X"F0",X"36",X"08",
		X"C3",X"85",X"24",X"3A",X"01",X"F0",X"C6",X"02",X"32",X"01",X"F0",X"FE",X"D0",X"C2",X"85",X"24",
		X"21",X"58",X"F0",X"36",X"09",X"FD",X"21",X"68",X"F8",X"FD",X"36",X"00",X"00",X"DD",X"36",X"04",
		X"FE",X"C3",X"85",X"24",X"DD",X"7E",X"07",X"D6",X"04",X"DD",X"77",X"07",X"CD",X"F3",X"43",X"DD",
		X"46",X"05",X"FD",X"21",X"5B",X"F2",X"CD",X"62",X"45",X"38",X"11",X"DD",X"36",X"0C",X"04",X"79",
		X"B7",X"3E",X"02",X"28",X"02",X"ED",X"44",X"DD",X"77",X"04",X"18",X"0C",X"21",X"58",X"F0",X"36",
		X"0A",X"DD",X"71",X"09",X"21",X"AF",X"F0",X"71",X"DD",X"7E",X"05",X"DD",X"86",X"04",X"DD",X"77",
		X"05",X"C3",X"85",X"24",X"DD",X"36",X"01",X"80",X"DD",X"7E",X"02",X"D6",X"16",X"FE",X"01",X"38",
		X"0B",X"28",X"12",X"21",X"FE",X"F0",X"36",X"03",X"3E",X"80",X"18",X"10",X"21",X"D2",X"F0",X"36",
		X"40",X"3E",X"08",X"18",X"07",X"21",X"D4",X"F0",X"36",X"03",X"3E",X"02",X"21",X"12",X"F0",X"B6",
		X"77",X"3A",X"5E",X"F0",X"B7",X"20",X"04",X"7E",X"EE",X"04",X"77",X"3E",X"04",X"32",X"5C",X"F0",
		X"DD",X"36",X"02",X"15",X"DD",X"36",X"06",X"29",X"DD",X"36",X"03",X"04",X"DD",X"36",X"0B",X"06",
		X"AF",X"32",X"5D",X"F0",X"32",X"58",X"F0",X"32",X"60",X"F0",X"32",X"03",X"F0",X"32",X"7F",X"F0",
		X"32",X"80",X"F0",X"3C",X"32",X"09",X"F4",X"3A",X"83",X"F0",X"EE",X"10",X"32",X"83",X"F0",X"21",
		X"06",X"F0",X"36",X"02",X"3A",X"7B",X"F3",X"B7",X"28",X"05",X"21",X"7A",X"F3",X"36",X"01",X"3A",
		X"33",X"F0",X"FE",X"03",X"C0",X"3A",X"34",X"F0",X"32",X"33",X"F0",X"C9",X"3A",X"01",X"F4",X"B7",
		X"C0",X"21",X"83",X"F0",X"46",X"DB",X"00",X"E6",X"10",X"77",X"23",X"70",X"3A",X"03",X"F0",X"47",
		X"E6",X"BB",X"28",X"14",X"2A",X"81",X"F0",X"3A",X"24",X"F0",X"B7",X"CA",X"E0",X"28",X"AF",X"32",
		X"24",X"F0",X"32",X"FC",X"F8",X"C3",X"E0",X"28",X"78",X"E6",X"40",X"28",X"13",X"2A",X"81",X"F0",
		X"7C",X"FE",X"04",X"DA",X"CB",X"28",X"7D",X"D6",X"04",X"30",X"01",X"25",X"6F",X"C3",X"CB",X"28",
		X"3A",X"7E",X"F0",X"47",X"B7",X"28",X"17",X"3A",X"7A",X"F3",X"FE",X"02",X"20",X"10",X"3D",X"32",
		X"7A",X"F3",X"32",X"8A",X"F3",X"AF",X"21",X"8B",X"F3",X"77",X"23",X"77",X"23",X"77",X"3A",X"83",
		X"F0",X"FE",X"10",X"28",X"28",X"3A",X"1A",X"F0",X"B7",X"20",X"11",X"3A",X"84",X"F0",X"FE",X"10",
		X"28",X"0A",X"3A",X"80",X"F0",X"FE",X"08",X"F2",X"5D",X"28",X"18",X"08",X"3A",X"80",X"F0",X"FE",
		X"12",X"F2",X"5D",X"28",X"3E",X"01",X"32",X"1A",X"F0",X"06",X"00",X"18",X"04",X"AF",X"32",X"1A",
		X"F0",X"ED",X"5B",X"7F",X"F0",X"7B",X"2F",X"6F",X"7A",X"2F",X"67",X"23",X"0E",X"00",X"09",X"0E",
		X"04",X"78",X"B7",X"28",X"1A",X"3A",X"83",X"F0",X"FE",X"10",X"28",X"13",X"78",X"FE",X"1F",X"38",
		X"0D",X"3A",X"1A",X"F0",X"B7",X"20",X"07",X"CD",X"6C",X"29",X"0D",X"41",X"18",X"0F",X"0C",X"41",
		X"3A",X"24",X"F0",X"B7",X"28",X"07",X"AF",X"32",X"24",X"F0",X"32",X"FC",X"F8",X"CB",X"2C",X"CB",
		X"1D",X"10",X"FA",X"19",X"3A",X"84",X"F0",X"47",X"3A",X"83",X"F0",X"B8",X"28",X"0B",X"FE",X"00",
		X"28",X"03",X"29",X"18",X"04",X"CB",X"2C",X"CB",X"1D",X"22",X"7F",X"F0",X"CB",X"2C",X"CB",X"1D",
		X"3A",X"83",X"F0",X"FE",X"00",X"28",X"04",X"CB",X"2C",X"CB",X"1D",X"22",X"81",X"F0",X"7C",X"B7",
		X"20",X"0E",X"3A",X"19",X"F0",X"47",X"3A",X"18",X"F0",X"B0",X"28",X"04",X"24",X"22",X"81",X"F0",
		X"3A",X"09",X"F4",X"FE",X"01",X"D8",X"20",X"72",X"3A",X"03",X"F0",X"E6",X"81",X"C0",X"3A",X"83",
		X"F0",X"FE",X"10",X"7C",X"28",X"02",X"C6",X"0D",X"6F",X"CB",X"27",X"85",X"47",X"3A",X"15",X"F0",
		X"21",X"05",X"2A",X"B7",X"28",X"03",X"21",X"5F",X"2A",X"78",X"85",X"30",X"01",X"24",X"6F",X"E5",
		X"FD",X"E1",X"3A",X"06",X"F4",X"FD",X"BE",X"00",X"20",X"15",X"FE",X"1F",X"C8",X"3A",X"07",X"F4",
		X"FD",X"BE",X"01",X"20",X"07",X"3A",X"08",X"F4",X"FD",X"BE",X"02",X"C8",X"3A",X"06",X"F4",X"FE",
		X"1F",X"20",X"05",X"0E",X"20",X"CD",X"4E",X"3D",X"FD",X"7E",X"00",X"32",X"06",X"F4",X"FE",X"1F",
		X"20",X"05",X"4F",X"CD",X"4E",X"3D",X"C9",X"4F",X"FD",X"7E",X"01",X"32",X"07",X"F4",X"57",X"FD",
		X"7E",X"02",X"32",X"08",X"F4",X"5F",X"CD",X"8E",X"3D",X"C9",X"0E",X"43",X"3A",X"15",X"F0",X"B7",
		X"28",X"02",X"0E",X"4A",X"CD",X"4E",X"3D",X"AF",X"32",X"09",X"F4",X"C9",X"3A",X"D5",X"F0",X"B7",
		X"C0",X"3A",X"24",X"F0",X"FE",X"04",X"D0",X"E5",X"47",X"CB",X"27",X"80",X"21",X"97",X"29",X"85",
		X"30",X"01",X"24",X"6F",X"FD",X"21",X"FC",X"F8",X"E9",X"3A",X"82",X"F0",X"FE",X"0F",X"38",X"05",
		X"21",X"24",X"F0",X"36",X"03",X"E1",X"C9",X"C3",X"A3",X"29",X"C3",X"B2",X"29",X"C3",X"D1",X"29",
		X"C3",X"EE",X"29",X"21",X"56",X"F1",X"36",X"10",X"21",X"24",X"F0",X"34",X"FD",X"36",X"01",X"00",
		X"18",X"D7",X"3A",X"56",X"F1",X"3D",X"28",X"0E",X"32",X"56",X"F1",X"E6",X"04",X"28",X"02",X"3E",
		X"7B",X"FD",X"77",X"02",X"18",X"C3",X"21",X"56",X"F1",X"36",X"10",X"21",X"24",X"F0",X"34",X"18",
		X"B8",X"3A",X"56",X"F1",X"3D",X"28",X"0F",X"32",X"56",X"F1",X"E6",X"02",X"28",X"02",X"3E",X"7B",
		X"FD",X"77",X"02",X"C3",X"89",X"29",X"21",X"56",X"F1",X"36",X"10",X"C3",X"89",X"29",X"FD",X"36",
		X"00",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"00",X"FD",X"36",X"03",X"00",X"21",X"24",
		X"F0",X"34",X"C3",X"95",X"29",X"BC",X"CF",X"F0",X"BC",X"CF",X"A0",X"BC",X"CF",X"50",X"BC",X"CF",
		X"00",X"BE",X"CE",X"C0",X"BE",X"CE",X"80",X"BE",X"CE",X"40",X"BE",X"CE",X"00",X"BE",X"CD",X"C0",
		X"BE",X"CD",X"C0",X"BE",X"CD",X"C0",X"BE",X"CD",X"C0",X"BE",X"CD",X"C0",X"1F",X"00",X"00",X"1F",
		X"00",X"00",X"1F",X"00",X"00",X"C0",X"CE",X"40",X"C0",X"CE",X"00",X"C0",X"CD",X"C0",X"C0",X"CD",
		X"80",X"C0",X"CD",X"40",X"C0",X"CD",X"00",X"C0",X"CC",X"C0",X"C0",X"CC",X"80",X"C2",X"CC",X"40",
		X"C2",X"CC",X"00",X"C2",X"CB",X"C0",X"C2",X"CB",X"80",X"C2",X"CB",X"40",X"C2",X"CB",X"00",X"C6",
		X"CF",X"F0",X"C6",X"CF",X"A0",X"C6",X"CF",X"50",X"C6",X"CF",X"00",X"C7",X"CE",X"C0",X"C7",X"CE",
		X"80",X"C7",X"CE",X"40",X"C7",X"CE",X"00",X"C7",X"CD",X"C0",X"C7",X"CD",X"C0",X"C7",X"CD",X"C0",
		X"C7",X"CD",X"C0",X"C7",X"CD",X"C0",X"1F",X"00",X"00",X"1F",X"00",X"00",X"1F",X"00",X"00",X"C8",
		X"CE",X"40",X"C8",X"CE",X"00",X"C8",X"CD",X"C0",X"C8",X"CD",X"80",X"C8",X"CD",X"40",X"C8",X"CD",
		X"00",X"C8",X"CC",X"C0",X"C8",X"CC",X"80",X"C9",X"CC",X"40",X"C9",X"CC",X"00",X"C9",X"CB",X"C0",
		X"C9",X"CB",X"80",X"C9",X"CB",X"40",X"C9",X"CB",X"00",X"3A",X"B8",X"F0",X"B7",X"C4",X"CC",X"2F",
		X"2A",X"81",X"F0",X"ED",X"5B",X"85",X"F0",X"19",X"7C",X"26",X"00",X"22",X"85",X"F0",X"B7",X"C8",
		X"F3",X"47",X"3A",X"0A",X"F0",X"B7",X"28",X"74",X"57",X"21",X"0D",X"F0",X"3A",X"A1",X"F0",X"CB",
		X"7A",X"20",X"27",X"B7",X"20",X"03",X"3C",X"18",X"15",X"CB",X"7F",X"28",X"11",X"ED",X"44",X"4F",
		X"3A",X"00",X"F0",X"81",X"FE",X"F0",X"38",X"02",X"3E",X"F0",X"32",X"00",X"F0",X"AF",X"4F",X"86",
		X"30",X"2D",X"3E",X"FF",X"96",X"4F",X"3E",X"FF",X"18",X"25",X"B7",X"28",X"3F",X"CB",X"7F",X"20",
		X"15",X"ED",X"44",X"4F",X"3A",X"00",X"F0",X"81",X"FE",X"10",X"30",X"02",X"3E",X"10",X"32",X"00",
		X"F0",X"0E",X"00",X"7E",X"18",X"09",X"4F",X"86",X"38",X"05",X"7E",X"ED",X"44",X"4F",X"AF",X"77",
		X"79",X"32",X"0C",X"F0",X"B7",X"28",X"15",X"3A",X"00",X"F0",X"82",X"CB",X"7A",X"20",X"06",X"FE",
		X"80",X"30",X"09",X"18",X"04",X"FE",X"80",X"38",X"03",X"32",X"00",X"F0",X"CD",X"CB",X"2B",X"CD",
		X"40",X"2C",X"2A",X"91",X"F0",X"2B",X"7C",X"E6",X"07",X"67",X"22",X"91",X"F0",X"21",X"87",X"F0",
		X"34",X"7E",X"FE",X"08",X"20",X"2F",X"3A",X"15",X"F0",X"B7",X"28",X"06",X"21",X"0B",X"F0",X"34",
		X"18",X"48",X"3A",X"0A",X"F0",X"B7",X"20",X"42",X"3A",X"14",X"F0",X"B7",X"20",X"3C",X"21",X"CE",
		X"F0",X"35",X"20",X"36",X"21",X"CF",X"F0",X"36",X"01",X"CD",X"E7",X"3C",X"E6",X"3F",X"C6",X"40",
		X"32",X"CE",X"F0",X"18",X"25",X"FE",X"10",X"20",X"21",X"36",X"00",X"3A",X"88",X"F0",X"B7",X"20",
		X"0E",X"3A",X"15",X"F0",X"B7",X"28",X"05",X"CD",X"E1",X"2E",X"18",X"03",X"CD",X"01",X"2E",X"DD",
		X"2A",X"93",X"F0",X"CD",X"41",X"46",X"DD",X"22",X"93",X"F0",X"10",X"96",X"3A",X"CF",X"F0",X"B7",
		X"28",X"07",X"CD",X"E4",X"3F",X"AF",X"32",X"CF",X"F0",X"FB",X"C9",X"21",X"AD",X"F0",X"48",X"11",
		X"04",X"00",X"DD",X"21",X"04",X"F8",X"06",X"14",X"3A",X"15",X"F0",X"B7",X"28",X"02",X"06",X"11",
		X"DD",X"7E",X"00",X"B7",X"28",X"54",X"3A",X"0C",X"F0",X"B7",X"28",X"0E",X"DD",X"86",X"00",X"FE",
		X"05",X"38",X"14",X"FE",X"F8",X"30",X"10",X"DD",X"77",X"00",X"DD",X"7E",X"03",X"81",X"38",X"07",
		X"DD",X"77",X"03",X"FE",X"F8",X"38",X"33",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"00",X"35",
		X"3A",X"EF",X"F0",X"B7",X"28",X"24",X"3A",X"FB",X"F0",X"B7",X"28",X"1E",X"FD",X"2A",X"FA",X"F0",
		X"FD",X"7E",X"02",X"DD",X"BE",X"02",X"20",X"12",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"20",X"0A",
		X"32",X"FB",X"F0",X"32",X"F5",X"F0",X"3C",X"32",X"F6",X"F0",X"DD",X"19",X"10",X"A2",X"41",X"C9",
		X"3A",X"9E",X"F0",X"FE",X"02",X"D8",X"48",X"06",X"03",X"28",X"02",X"06",X"06",X"DD",X"21",X"A8",
		X"F9",X"26",X"00",X"DD",X"7E",X"00",X"B7",X"28",X"44",X"3A",X"0C",X"F0",X"B7",X"28",X"0E",X"DD",
		X"86",X"00",X"FE",X"05",X"38",X"11",X"FE",X"F8",X"30",X"0D",X"DD",X"77",X"00",X"DD",X"7E",X"03",
		X"81",X"38",X"04",X"FE",X"F8",X"38",X"0E",X"DD",X"36",X"00",X"00",X"DD",X"36",X"02",X"19",X"DD",
		X"36",X"01",X"00",X"18",X"18",X"6F",X"3A",X"15",X"F0",X"57",X"3A",X"06",X"F0",X"BA",X"20",X"09",
		X"3A",X"01",X"F0",X"DD",X"BE",X"03",X"DC",X"AD",X"2C",X"DD",X"75",X"03",X"24",X"11",X"04",X"00",
		X"DD",X"19",X"10",X"AF",X"7C",X"B7",X"20",X"03",X"32",X"9E",X"F0",X"41",X"C9",X"E5",X"3A",X"17",
		X"F0",X"B7",X"CA",X"BE",X"2D",X"C5",X"DD",X"E5",X"21",X"A6",X"F0",X"36",X"11",X"AF",X"32",X"17",
		X"F0",X"32",X"45",X"F0",X"3A",X"16",X"F0",X"B7",X"28",X"63",X"CD",X"01",X"56",X"AF",X"32",X"46",
		X"F0",X"32",X"18",X"F0",X"32",X"FC",X"F8",X"32",X"0B",X"F0",X"32",X"22",X"F0",X"32",X"0C",X"F0",
		X"32",X"0D",X"F0",X"32",X"56",X"F0",X"32",X"42",X"F0",X"32",X"57",X"F0",X"32",X"60",X"F0",X"32",
		X"5E",X"F0",X"32",X"60",X"F8",X"32",X"64",X"F8",X"3C",X"32",X"15",X"F0",X"32",X"0A",X"F0",X"3A",
		X"03",X"F0",X"F6",X"40",X"32",X"03",X"F0",X"21",X"04",X"F0",X"36",X"1C",X"21",X"02",X"F0",X"36",
		X"08",X"3A",X"12",X"F0",X"E6",X"8B",X"32",X"12",X"F0",X"21",X"82",X"F0",X"7E",X"FE",X"0C",X"38",
		X"04",X"36",X"0C",X"18",X"4C",X"FE",X"04",X"30",X"48",X"36",X"04",X"18",X"44",X"32",X"0C",X"F0",
		X"32",X"19",X"F0",X"32",X"81",X"F0",X"32",X"82",X"F0",X"32",X"7F",X"F0",X"32",X"80",X"F0",X"32",
		X"00",X"F0",X"DD",X"21",X"6C",X"F8",X"DD",X"77",X"00",X"DD",X"77",X"04",X"32",X"B9",X"F0",X"3D",
		X"32",X"0A",X"F0",X"32",X"0D",X"F0",X"3A",X"03",X"F0",X"F6",X"10",X"32",X"03",X"F0",X"21",X"09",
		X"F4",X"36",X"02",X"21",X"90",X"F3",X"34",X"21",X"B8",X"F0",X"36",X"01",X"21",X"04",X"F0",X"36",
		X"14",X"DD",X"21",X"48",X"F8",X"11",X"04",X"00",X"06",X"06",X"AF",X"DD",X"77",X"00",X"DD",X"19",
		X"10",X"F9",X"3A",X"A0",X"F0",X"57",X"AF",X"32",X"A0",X"F0",X"DD",X"21",X"8B",X"F2",X"1E",X"00",
		X"01",X"23",X"00",X"DD",X"7E",X"01",X"E6",X"80",X"28",X"17",X"DD",X"7E",X"05",X"B7",X"20",X"05",
		X"CD",X"32",X"3F",X"18",X"0C",X"7A",X"B7",X"28",X"08",X"DD",X"36",X"03",X"01",X"DD",X"36",X"0B",
		X"01",X"DD",X"09",X"1C",X"7B",X"FE",X"06",X"20",X"DA",X"DD",X"E1",X"C1",X"E1",X"C9",X"21",X"16",
		X"F0",X"3A",X"15",X"F0",X"BE",X"28",X"1E",X"B7",X"20",X"0F",X"21",X"02",X"F0",X"36",X"11",X"3A",
		X"03",X"F0",X"F6",X"40",X"32",X"03",X"F0",X"18",X"0C",X"AF",X"32",X"00",X"F0",X"3A",X"03",X"F0",
		X"F6",X"10",X"32",X"03",X"F0",X"E1",X"C9",X"7D",X"C6",X"10",X"6F",X"D0",X"7C",X"3C",X"E6",X"E3",
		X"67",X"C9",X"7D",X"D6",X"10",X"6F",X"D0",X"7C",X"3D",X"FE",X"E0",X"30",X"02",X"3E",X"E3",X"67",
		X"C9",X"3A",X"18",X"F0",X"FE",X"01",X"D8",X"C5",X"20",X"59",X"3D",X"32",X"17",X"F0",X"0E",X"10",
		X"06",X"C0",X"CD",X"21",X"72",X"7E",X"FE",X"42",X"28",X"02",X"C1",X"C9",X"23",X"22",X"9B",X"F0",
		X"06",X"07",X"36",X"02",X"CD",X"E7",X"2D",X"10",X"F9",X"36",X"6F",X"CD",X"E7",X"2D",X"36",X"D3",
		X"CD",X"E7",X"2D",X"36",X"7B",X"CD",X"E7",X"2D",X"36",X"D0",X"06",X"31",X"CD",X"E7",X"2D",X"36",
		X"AF",X"10",X"F9",X"CD",X"E7",X"2D",X"36",X"E8",X"CD",X"E7",X"2D",X"36",X"02",X"CD",X"E7",X"2D",
		X"36",X"01",X"CD",X"E7",X"2D",X"36",X"40",X"21",X"18",X"F0",X"36",X"02",X"3E",X"01",X"32",X"16",
		X"F0",X"C1",X"C9",X"FE",X"03",X"28",X"06",X"3C",X"32",X"18",X"F0",X"C1",X"C9",X"2A",X"9B",X"F0",
		X"7C",X"F6",X"04",X"67",X"7D",X"E6",X"F0",X"6F",X"11",X"0E",X"1C",X"19",X"22",X"97",X"F0",X"21",
		X"18",X"F0",X"34",X"AF",X"32",X"09",X"F0",X"32",X"8A",X"F0",X"32",X"8B",X"F0",X"32",X"89",X"F0",
		X"32",X"8F",X"F0",X"32",X"90",X"F0",X"3C",X"32",X"17",X"F0",X"32",X"A3",X"F0",X"DD",X"21",X"E9",
		X"BE",X"DD",X"22",X"99",X"F0",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"22",X"3C",X"F0",X"DD",X"6E",
		X"04",X"DD",X"66",X"05",X"5E",X"23",X"56",X"ED",X"53",X"95",X"F0",X"23",X"7E",X"DD",X"21",X"61",
		X"F0",X"DD",X"77",X"01",X"DD",X"36",X"02",X"40",X"11",X"03",X"00",X"ED",X"53",X"7C",X"F0",X"23",
		X"23",X"E5",X"DD",X"E1",X"06",X"7E",X"CD",X"41",X"46",X"10",X"FB",X"DD",X"22",X"93",X"F0",X"C1",
		X"C9",X"3A",X"19",X"F0",X"FE",X"01",X"D8",X"C5",X"20",X"67",X"3D",X"32",X"17",X"F0",X"0E",X"F0",
		X"06",X"C0",X"CD",X"21",X"72",X"7E",X"FE",X"1F",X"28",X"02",X"C1",X"C9",X"7C",X"E6",X"E3",X"67",
		X"7D",X"F6",X"0F",X"6F",X"CD",X"F2",X"2D",X"22",X"9B",X"F0",X"06",X"0C",X"36",X"02",X"CD",X"F2",
		X"2D",X"10",X"F9",X"36",X"85",X"CD",X"F2",X"2D",X"36",X"82",X"CD",X"F2",X"2D",X"36",X"38",X"CD",
		X"F2",X"2D",X"36",X"3E",X"CD",X"F2",X"2D",X"36",X"04",X"CD",X"F2",X"2D",X"36",X"33",X"CD",X"F2",
		X"2D",X"36",X"30",X"CD",X"F2",X"2D",X"36",X"34",X"CD",X"F2",X"2D",X"36",X"31",X"06",X"1B",X"CD",
		X"F2",X"2D",X"36",X"02",X"10",X"F9",X"21",X"19",X"F0",X"36",X"02",X"AF",X"32",X"16",X"F0",X"C1",
		X"C9",X"FE",X"03",X"28",X"06",X"3C",X"32",X"19",X"F0",X"C1",X"C9",X"2A",X"9B",X"F0",X"7D",X"E6",
		X"F0",X"6F",X"11",X"0E",X"20",X"19",X"22",X"97",X"F0",X"21",X"19",X"F0",X"34",X"AF",X"32",X"09",
		X"F0",X"32",X"8A",X"F0",X"32",X"8B",X"F0",X"32",X"89",X"F0",X"32",X"8F",X"F0",X"32",X"90",X"F0",
		X"3C",X"32",X"17",X"F0",X"DD",X"21",X"41",X"BF",X"DD",X"22",X"99",X"F0",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"22",X"3C",X"F0",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"5E",X"23",X"56",X"ED",X"53",
		X"95",X"F0",X"23",X"7E",X"DD",X"21",X"61",X"F0",X"DD",X"77",X"01",X"DD",X"36",X"02",X"40",X"11",
		X"03",X"00",X"ED",X"53",X"7C",X"F0",X"23",X"23",X"E5",X"DD",X"E1",X"06",X"7E",X"CD",X"41",X"46",
		X"10",X"FB",X"DD",X"22",X"93",X"F0",X"AF",X"32",X"33",X"F0",X"C1",X"C9",X"3A",X"B9",X"F0",X"B7",
		X"28",X"04",X"DD",X"2A",X"B2",X"F0",X"47",X"CB",X"27",X"80",X"21",X"10",X"30",X"85",X"30",X"01",
		X"24",X"6F",X"E9",X"21",X"B9",X"F0",X"34",X"DD",X"7E",X"03",X"32",X"82",X"F0",X"DD",X"7E",X"04",
		X"ED",X"44",X"32",X"A1",X"F0",X"DD",X"35",X"0C",X"C0",X"DD",X"36",X"0C",X"06",X"DD",X"7E",X"06",
		X"06",X"29",X"B8",X"20",X"02",X"06",X"D3",X"DD",X"70",X"06",X"C9",X"21",X"B9",X"F0",X"34",X"C9",
		X"C3",X"2E",X"30",X"C3",X"B8",X"30",X"C3",X"CD",X"30",X"C3",X"E9",X"30",X"C3",X"08",X"31",X"C3",
		X"38",X"31",X"C3",X"74",X"31",X"C3",X"82",X"31",X"C3",X"95",X"31",X"C3",X"BB",X"31",X"DD",X"21",
		X"8B",X"F2",X"06",X"06",X"11",X"23",X"00",X"DD",X"7E",X"01",X"B7",X"28",X"0A",X"DD",X"19",X"10",
		X"F6",X"DD",X"21",X"8B",X"F2",X"18",X"04",X"21",X"32",X"F0",X"34",X"DD",X"22",X"B2",X"F0",X"FD",
		X"2A",X"B6",X"F0",X"FD",X"7E",X"00",X"DD",X"77",X"05",X"FD",X"7E",X"03",X"DD",X"77",X"07",X"DD",
		X"36",X"08",X"00",X"DD",X"36",X"02",X"15",X"DD",X"36",X"06",X"29",X"3A",X"E6",X"BA",X"DD",X"77",
		X"0E",X"3A",X"EF",X"BA",X"DD",X"77",X"0F",X"DD",X"36",X"01",X"01",X"DD",X"36",X"0B",X"06",X"AF",
		X"DD",X"77",X"1F",X"DD",X"77",X"0A",X"DD",X"77",X"1E",X"DD",X"77",X"04",X"DD",X"36",X"03",X"03",
		X"DD",X"36",X"0D",X"15",X"DD",X"36",X"0C",X"01",X"FD",X"77",X"00",X"FD",X"2A",X"B4",X"F0",X"FD",
		X"46",X"02",X"DD",X"70",X"1D",X"FD",X"77",X"00",X"3A",X"AD",X"F0",X"D6",X"02",X"32",X"AD",X"F0",
		X"21",X"09",X"F4",X"36",X"02",X"C3",X"E3",X"2F",X"DD",X"35",X"0D",X"C2",X"F5",X"2F",X"DD",X"36",
		X"0D",X"30",X"DD",X"36",X"03",X"04",X"DD",X"36",X"04",X"01",X"C3",X"E3",X"2F",X"DD",X"35",X"0D",
		X"28",X"10",X"21",X"09",X"F4",X"36",X"02",X"DD",X"7E",X"04",X"EE",X"01",X"DD",X"77",X"04",X"C3",
		X"ED",X"2F",X"DD",X"36",X"04",X"01",X"C3",X"E3",X"2F",X"3A",X"0A",X"F0",X"B7",X"C2",X"F5",X"2F",
		X"32",X"15",X"F0",X"32",X"81",X"F0",X"32",X"82",X"F0",X"32",X"85",X"F0",X"32",X"86",X"F0",X"32",
		X"A1",X"F0",X"CD",X"F5",X"2F",X"C3",X"0B",X"30",X"DD",X"7E",X"07",X"D6",X"03",X"DD",X"77",X"07",
		X"DD",X"7E",X"05",X"3C",X"DD",X"77",X"05",X"FE",X"E5",X"C2",X"F5",X"2F",X"DD",X"36",X"04",X"00",
		X"DD",X"7E",X"07",X"FE",X"A0",X"3E",X"00",X"28",X"06",X"3E",X"02",X"38",X"02",X"ED",X"44",X"DD",
		X"77",X"03",X"CD",X"F5",X"2F",X"C3",X"0B",X"30",X"DD",X"7E",X"07",X"DD",X"86",X"03",X"DD",X"77",
		X"07",X"FE",X"A0",X"DA",X"F5",X"2F",X"DD",X"36",X"07",X"A0",X"DD",X"36",X"06",X"29",X"21",X"00",
		X"F0",X"DD",X"7E",X"05",X"77",X"32",X"07",X"F0",X"23",X"36",X"AC",X"23",X"36",X"08",X"DD",X"36",
		X"0D",X"10",X"FD",X"21",X"68",X"F8",X"FD",X"77",X"00",X"FD",X"36",X"02",X"2B",X"FD",X"36",X"03",
		X"B0",X"C3",X"0B",X"30",X"FD",X"21",X"68",X"F8",X"FD",X"34",X"03",X"DD",X"35",X"0D",X"C0",X"C3",
		X"0B",X"30",X"3A",X"01",X"F0",X"C6",X"02",X"32",X"01",X"F0",X"FE",X"D0",X"C0",X"21",X"68",X"F8",
		X"36",X"00",X"C3",X"0B",X"30",X"DD",X"7E",X"07",X"D6",X"04",X"DD",X"77",X"07",X"CD",X"F3",X"43",
		X"DD",X"7E",X"05",X"D6",X"02",X"DD",X"77",X"05",X"47",X"FD",X"21",X"5B",X"F2",X"CD",X"62",X"45",
		X"D0",X"DD",X"71",X"09",X"21",X"AF",X"F0",X"71",X"C3",X"0B",X"30",X"DD",X"36",X"01",X"80",X"DD",
		X"36",X"04",X"FE",X"DD",X"36",X"0C",X"04",X"DD",X"36",X"03",X"04",X"DD",X"36",X"0D",X"04",X"21",
		X"06",X"F0",X"36",X"02",X"21",X"05",X"F0",X"36",X"04",X"AF",X"32",X"03",X"F0",X"32",X"B9",X"F0",
		X"32",X"B8",X"F0",X"3A",X"8E",X"F3",X"FE",X"07",X"38",X"02",X"3E",X"07",X"2A",X"30",X"F0",X"85",
		X"30",X"01",X"24",X"6F",X"7E",X"32",X"33",X"F0",X"3E",X"02",X"32",X"35",X"F0",X"DD",X"7E",X"1D",
		X"FE",X"6A",X"20",X"09",X"21",X"D2",X"F0",X"36",X"40",X"3E",X"08",X"18",X"14",X"FE",X"6B",X"20",
		X"09",X"21",X"D4",X"F0",X"36",X"03",X"3E",X"02",X"18",X"07",X"21",X"FE",X"F0",X"36",X"03",X"3E",
		X"80",X"21",X"12",X"F0",X"B6",X"77",X"21",X"09",X"F4",X"36",X"01",X"3A",X"83",X"F0",X"EE",X"10",
		X"32",X"83",X"F0",X"C9",X"CD",X"41",X"32",X"CD",X"ED",X"36",X"CD",X"81",X"38",X"CD",X"2C",X"39",
		X"C9",X"AF",X"32",X"AE",X"F0",X"0E",X"00",X"FD",X"21",X"04",X"F8",X"21",X"41",X"F1",X"22",X"57",
		X"F1",X"FD",X"7E",X"00",X"B7",X"CA",X"53",X"36",X"7E",X"E6",X"0F",X"47",X"CA",X"40",X"36",X"FE",
		X"07",X"20",X"19",X"7E",X"D6",X"10",X"77",X"FE",X"07",X"20",X"0E",X"36",X"67",X"26",X"75",X"FD",
		X"7E",X"02",X"BC",X"20",X"01",X"24",X"FD",X"74",X"02",X"78",X"18",X"23",X"FE",X"08",X"20",X"1F",
		X"3A",X"AE",X"F0",X"3C",X"32",X"AE",X"F0",X"7E",X"D6",X"10",X"77",X"FE",X"08",X"20",X"0F",X"36",
		X"28",X"FD",X"7E",X"02",X"3C",X"FE",X"A0",X"38",X"02",X"3E",X"9C",X"FD",X"77",X"02",X"78",X"CB",
		X"27",X"CB",X"27",X"21",X"4D",X"BB",X"85",X"30",X"01",X"24",X"6F",X"E5",X"DD",X"E1",X"FD",X"7E",
		X"00",X"DD",X"86",X"00",X"57",X"FD",X"7E",X"03",X"DD",X"86",X"02",X"5F",X"3A",X"03",X"F0",X"E6",
		X"50",X"C2",X"22",X"34",X"7B",X"21",X"01",X"F0",X"DD",X"86",X"03",X"BE",X"DA",X"22",X"34",X"3A",
		X"04",X"F0",X"86",X"BB",X"DA",X"22",X"34",X"21",X"00",X"F0",X"7A",X"DD",X"86",X"01",X"BE",X"DA",
		X"22",X"34",X"7E",X"C6",X"10",X"BA",X"DA",X"22",X"34",X"78",X"FE",X"03",X"30",X"6B",X"FE",X"02",
		X"28",X"0C",X"1E",X"20",X"7E",X"BA",X"30",X"19",X"1E",X"00",X"C6",X"10",X"18",X"15",X"1E",X"00",
		X"7A",X"DD",X"86",X"01",X"57",X"7E",X"C6",X"10",X"BA",X"38",X"08",X"1E",X"20",X"D6",X"20",X"18",
		X"02",X"D6",X"10",X"FD",X"77",X"00",X"FD",X"7E",X"03",X"D6",X"08",X"FD",X"77",X"03",X"FD",X"73",
		X"01",X"FD",X"36",X"02",X"13",X"2A",X"57",X"F1",X"36",X"50",X"3A",X"02",X"F0",X"FE",X"08",X"C2",
		X"53",X"36",X"3A",X"03",X"F0",X"F6",X"04",X"32",X"03",X"F0",X"CD",X"E7",X"3C",X"5F",X"3E",X"02",
		X"16",X"07",X"CB",X"43",X"28",X"04",X"ED",X"44",X"16",X"00",X"32",X"A1",X"F0",X"21",X"02",X"F0",
		X"72",X"21",X"27",X"F0",X"36",X"06",X"C3",X"53",X"36",X"CA",X"53",X"36",X"FE",X"06",X"28",X"36",
		X"FE",X"05",X"CA",X"E9",X"33",X"FE",X"07",X"20",X"11",X"3A",X"82",X"F0",X"FE",X"05",X"DA",X"53",
		X"36",X"FD",X"36",X"02",X"39",X"2A",X"57",X"F1",X"36",X"50",X"C5",X"0E",X"13",X"CD",X"4E",X"3D",
		X"FD",X"E5",X"CD",X"CB",X"7D",X"FD",X"E1",X"C1",X"3A",X"56",X"F0",X"B7",X"C2",X"53",X"36",X"3C",
		X"32",X"56",X"F0",X"C3",X"53",X"36",X"3A",X"A1",X"F0",X"ED",X"44",X"20",X"0C",X"3A",X"00",X"F0",
		X"FD",X"BE",X"00",X"3E",X"08",X"38",X"02",X"ED",X"44",X"FD",X"86",X"00",X"FD",X"77",X"00",X"3A",
		X"15",X"F0",X"B7",X"28",X"34",X"FD",X"7E",X"02",X"FE",X"BB",X"28",X"04",X"FE",X"BF",X"20",X"06",
		X"DD",X"2A",X"2C",X"F0",X"18",X"0C",X"FE",X"BC",X"28",X"04",X"FE",X"C0",X"20",X"1B",X"DD",X"2A",
		X"2A",X"F0",X"FD",X"7E",X"00",X"DD",X"96",X"00",X"30",X"02",X"ED",X"44",X"FE",X"09",X"30",X"09",
		X"FD",X"7E",X"00",X"DD",X"77",X"00",X"CD",X"6F",X"36",X"3A",X"82",X"F0",X"FE",X"07",X"38",X"23",
		X"3A",X"03",X"F0",X"F6",X"02",X"32",X"03",X"F0",X"21",X"A1",X"F0",X"3A",X"00",X"F0",X"FE",X"80",
		X"3E",X"02",X"30",X"02",X"ED",X"44",X"77",X"3A",X"06",X"F0",X"FE",X"02",X"C2",X"13",X"34",X"AF",
		X"32",X"06",X"F0",X"C5",X"0E",X"12",X"CD",X"4E",X"3D",X"C1",X"3E",X"01",X"32",X"09",X"F0",X"C3",
		X"53",X"36",X"C5",X"FD",X"E5",X"0E",X"00",X"FD",X"21",X"8B",X"F2",X"FD",X"7E",X"08",X"B7",X"C2",
		X"30",X"36",X"FD",X"7E",X"05",X"B7",X"CA",X"30",X"36",X"C6",X"10",X"BA",X"DA",X"30",X"36",X"7A",
		X"DD",X"86",X"01",X"FD",X"BE",X"05",X"DA",X"30",X"36",X"FD",X"7E",X"07",X"FD",X"86",X"0E",X"DA",
		X"30",X"36",X"BB",X"DA",X"30",X"36",X"7B",X"DD",X"86",X"03",X"DA",X"30",X"36",X"FD",X"BE",X"07",
		X"DA",X"30",X"36",X"FD",X"6E",X"05",X"FD",X"22",X"3A",X"F0",X"FD",X"E1",X"78",X"FE",X"03",X"D2",
		X"49",X"35",X"FE",X"02",X"28",X"0C",X"1E",X"20",X"7D",X"BA",X"30",X"1D",X"1E",X"00",X"C6",X"14",
		X"18",X"19",X"1E",X"00",X"7A",X"DD",X"86",X"01",X"57",X"7D",X"C6",X"10",X"BA",X"38",X"06",X"1E",
		X"20",X"D6",X"24",X"18",X"06",X"C6",X"04",X"18",X"02",X"D6",X"14",X"FD",X"77",X"00",X"FD",X"7E",
		X"03",X"D6",X"08",X"FD",X"77",X"03",X"FD",X"73",X"01",X"FD",X"36",X"02",X"13",X"2A",X"57",X"F1",
		X"36",X"50",X"DD",X"2A",X"3A",X"F0",X"DD",X"7E",X"0C",X"C6",X"03",X"DD",X"77",X"0C",X"18",X"6F",
		X"DD",X"7E",X"01",X"E6",X"04",X"28",X"08",X"DD",X"7E",X"0C",X"FE",X"60",X"D2",X"52",X"36",X"DD",
		X"36",X"0C",X"80",X"DD",X"36",X"21",X"00",X"DD",X"36",X"22",X"02",X"3A",X"15",X"F0",X"B7",X"20",
		X"1F",X"3A",X"82",X"F0",X"3D",X"DD",X"77",X"03",X"FE",X"08",X"30",X"14",X"3A",X"49",X"F0",X"B7",
		X"20",X"0E",X"21",X"45",X"F0",X"7E",X"B7",X"20",X"07",X"36",X"03",X"21",X"42",X"F0",X"36",X"01",
		X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"01",X"20",X"10",X"DD",X"7E",X"06",X"FE",X"7C",X"3E",X"00",
		X"28",X"02",X"C6",X"04",X"DD",X"77",X"16",X"18",X"16",X"FE",X"06",X"38",X"12",X"3A",X"12",X"F0",
		X"E6",X"FB",X"32",X"12",X"F0",X"AF",X"32",X"5C",X"F0",X"32",X"58",X"F0",X"32",X"5E",X"F0",X"DD",
		X"7E",X"01",X"F6",X"04",X"DD",X"77",X"01",X"DD",X"36",X"0D",X"10",X"3E",X"02",X"CB",X"41",X"28",
		X"02",X"ED",X"44",X"DD",X"77",X"04",X"C3",X"52",X"36",X"DD",X"2A",X"3A",X"F0",X"CA",X"C0",X"34",
		X"FE",X"06",X"28",X"5B",X"FE",X"04",X"28",X"36",X"FE",X"07",X"28",X"29",X"FE",X"08",X"DD",X"7E",
		X"02",X"20",X"11",X"67",X"DD",X"7E",X"01",X"E6",X"02",X"C2",X"52",X"36",X"7C",X"C5",X"CD",X"91",
		X"3E",X"C1",X"18",X"1A",X"E6",X"0F",X"FE",X"05",X"D2",X"52",X"36",X"DD",X"7E",X"01",X"F6",X"02",
		X"DD",X"77",X"01",X"18",X"B6",X"FD",X"36",X"02",X"39",X"2A",X"57",X"F1",X"36",X"50",X"DD",X"7E",
		X"02",X"E6",X"0F",X"FE",X"05",X"D2",X"52",X"36",X"DD",X"7E",X"01",X"E6",X"03",X"FE",X"03",X"28",
		X"9A",X"DD",X"7E",X"01",X"F6",X"03",X"DD",X"77",X"01",X"DD",X"36",X"1F",X"10",X"18",X"8C",X"C5",
		X"0E",X"12",X"CD",X"4E",X"3D",X"C1",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"05",X"30",X"08",X"DD",
		X"7E",X"01",X"F6",X"02",X"DD",X"77",X"01",X"DD",X"7E",X"05",X"FD",X"BE",X"00",X"3E",X"08",X"38",
		X"08",X"ED",X"44",X"DD",X"36",X"04",X"02",X"18",X"04",X"DD",X"36",X"04",X"FE",X"FD",X"86",X"00",
		X"FD",X"77",X"00",X"3A",X"15",X"F0",X"B7",X"28",X"3A",X"FD",X"7E",X"02",X"FE",X"BB",X"28",X"04",
		X"FE",X"BF",X"20",X"08",X"DD",X"E5",X"DD",X"2A",X"2C",X"F0",X"18",X"0E",X"FE",X"BC",X"28",X"04",
		X"FE",X"C0",X"20",X"1F",X"DD",X"E5",X"DD",X"2A",X"2A",X"F0",X"FD",X"7E",X"00",X"DD",X"96",X"00",
		X"30",X"02",X"ED",X"44",X"FE",X"09",X"30",X"09",X"FD",X"7E",X"00",X"DD",X"77",X"00",X"CD",X"6F",
		X"36",X"DD",X"E1",X"DD",X"7E",X"10",X"CB",X"27",X"FD",X"86",X"03",X"FD",X"77",X"03",X"18",X"22",
		X"D5",X"11",X"23",X"00",X"FD",X"19",X"D1",X"0C",X"79",X"FE",X"06",X"C2",X"2B",X"34",X"18",X"10",
		X"7E",X"D6",X"10",X"77",X"20",X"0D",X"FD",X"36",X"00",X"00",X"21",X"AD",X"F0",X"35",X"18",X"03",
		X"FD",X"E1",X"C1",X"0C",X"3A",X"15",X"F0",X"B7",X"3E",X"14",X"28",X"02",X"D6",X"03",X"B9",X"C8",
		X"11",X"04",X"00",X"FD",X"19",X"2A",X"57",X"F1",X"23",X"22",X"57",X"F1",X"C3",X"51",X"32",X"3A",
		X"B0",X"F0",X"B7",X"C0",X"FD",X"E5",X"DD",X"E5",X"C5",X"06",X"00",X"FD",X"2A",X"2C",X"F0",X"FD",
		X"4E",X"03",X"FD",X"21",X"5B",X"F2",X"CD",X"B5",X"41",X"2A",X"2A",X"F0",X"46",X"CD",X"62",X"45",
		X"47",X"3E",X"01",X"38",X"0F",X"16",X"02",X"79",X"B7",X"20",X"02",X"14",X"78",X"FE",X"0C",X"3E",
		X"00",X"30",X"01",X"82",X"57",X"FE",X"01",X"FD",X"2A",X"2A",X"F0",X"DD",X"2A",X"2C",X"F0",X"30",
		X"0E",X"FD",X"36",X"02",X"BF",X"DD",X"36",X"00",X"00",X"21",X"AD",X"F0",X"35",X"18",X"28",X"20",
		X"12",X"FD",X"36",X"00",X"00",X"DD",X"36",X"00",X"00",X"3A",X"AD",X"F0",X"D6",X"02",X"32",X"AD",
		X"F0",X"18",X"14",X"FD",X"36",X"02",X"BB",X"DD",X"36",X"02",X"BC",X"FE",X"02",X"20",X"08",X"FD",
		X"36",X"01",X"20",X"DD",X"36",X"01",X"20",X"C1",X"DD",X"E1",X"FD",X"E1",X"C9",X"3A",X"EF",X"F0",
		X"B7",X"C8",X"FE",X"02",X"CA",X"CC",X"37",X"3A",X"F4",X"F0",X"21",X"F7",X"F0",X"86",X"32",X"F4",
		X"F0",X"3A",X"82",X"F0",X"21",X"F6",X"F0",X"46",X"21",X"F8",X"F0",X"96",X"21",X"F5",X"F0",X"CB",
		X"7F",X"28",X"06",X"86",X"38",X"07",X"05",X"18",X"04",X"86",X"30",X"01",X"04",X"77",X"78",X"32",
		X"F6",X"F0",X"FD",X"21",X"C0",X"F9",X"21",X"F0",X"F0",X"35",X"28",X"15",X"B7",X"20",X"0D",X"3A",
		X"F4",X"F0",X"FD",X"77",X"00",X"3A",X"F5",X"F0",X"FD",X"77",X"03",X"C9",X"FD",X"36",X"00",X"00",
		X"C9",X"FD",X"36",X"00",X"00",X"36",X"04",X"21",X"EF",X"F0",X"34",X"0E",X"17",X"CD",X"4E",X"3D",
		X"21",X"F9",X"F0",X"36",X"38",X"78",X"B7",X"20",X"68",X"CD",X"B3",X"3D",X"FD",X"36",X"02",X"38",
		X"CD",X"E4",X"3D",X"36",X"04",X"22",X"59",X"F1",X"FD",X"22",X"FA",X"F0",X"3A",X"15",X"F0",X"B7",
		X"28",X"3B",X"3A",X"0A",X"F0",X"B7",X"28",X"04",X"3E",X"01",X"18",X"31",X"3A",X"19",X"F0",X"B7",
		X"20",X"F6",X"3A",X"82",X"F0",X"B7",X"28",X"F0",X"06",X"00",X"21",X"F5",X"F0",X"4E",X"FD",X"21",
		X"5B",X"F2",X"CD",X"B5",X"41",X"21",X"F4",X"F0",X"46",X"CD",X"62",X"45",X"47",X"3E",X"01",X"38",
		X"0C",X"79",X"B7",X"20",X"01",X"78",X"FE",X"0C",X"3E",X"00",X"30",X"01",X"3C",X"32",X"F1",X"F0",
		X"FD",X"2A",X"FA",X"F0",X"3A",X"F4",X"F0",X"FD",X"77",X"00",X"3A",X"F5",X"F0",X"FD",X"77",X"03",
		X"C9",X"AF",X"32",X"FB",X"F0",X"3A",X"15",X"F0",X"32",X"F1",X"F0",X"C9",X"21",X"F0",X"F0",X"35",
		X"20",X"56",X"36",X"04",X"21",X"F9",X"F0",X"7E",X"FE",X"38",X"20",X"0A",X"3A",X"F1",X"F0",X"B7",
		X"28",X"10",X"36",X"A2",X"18",X"2C",X"FE",X"3D",X"28",X"0B",X"FE",X"A6",X"20",X"04",X"36",X"00",
		X"18",X"03",X"34",X"18",X"1D",X"0E",X"18",X"CD",X"4E",X"3D",X"3A",X"FB",X"F0",X"B7",X"20",X"16",
		X"3A",X"F9",X"F0",X"B7",X"28",X"6A",X"3A",X"F6",X"F0",X"FE",X"FF",X"28",X"20",X"B7",X"28",X"1D",
		X"18",X"5E",X"3A",X"FB",X"F0",X"B7",X"28",X"15",X"FD",X"2A",X"FA",X"F0",X"7E",X"FD",X"77",X"02",
		X"B7",X"28",X"52",X"FE",X"3D",X"C0",X"18",X"43",X"3A",X"FB",X"F0",X"B7",X"C0",X"21",X"82",X"F0",
		X"3A",X"F5",X"F0",X"86",X"21",X"F6",X"F0",X"30",X"01",X"34",X"32",X"F5",X"F0",X"3A",X"F6",X"F0",
		X"B7",X"C0",X"CD",X"B3",X"3D",X"FD",X"22",X"FA",X"F0",X"CD",X"E4",X"3D",X"22",X"59",X"F1",X"3A",
		X"F4",X"F0",X"FD",X"77",X"00",X"3A",X"F5",X"F0",X"FD",X"77",X"03",X"3A",X"F9",X"F0",X"FD",X"77",
		X"02",X"B7",X"28",X"11",X"FE",X"3D",X"28",X"03",X"36",X"04",X"C9",X"2A",X"59",X"F1",X"36",X"05",
		X"AF",X"32",X"EF",X"F0",X"C9",X"AF",X"FD",X"77",X"00",X"32",X"EF",X"F0",X"2A",X"59",X"F1",X"77",
		X"C9",X"3A",X"BA",X"F0",X"B7",X"28",X"17",X"DD",X"2A",X"BD",X"F0",X"21",X"A8",X"38",X"3D",X"47",
		X"CB",X"27",X"80",X"85",X"30",X"01",X"24",X"6F",X"E9",X"21",X"BA",X"F0",X"34",X"C9",X"3A",X"BB",
		X"F0",X"B7",X"C8",X"3D",X"32",X"BB",X"F0",X"C9",X"C3",X"B1",X"38",X"C3",X"E5",X"38",X"C3",X"0E",
		X"39",X"21",X"BB",X"F0",X"35",X"28",X"0A",X"3A",X"BC",X"F0",X"DD",X"86",X"03",X"DD",X"77",X"03",
		X"C9",X"36",X"03",X"CD",X"B3",X"3D",X"FD",X"22",X"BF",X"F0",X"CD",X"E4",X"3D",X"36",X"97",X"DD",
		X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"FD",X"36",X"02",X"A3",X"FD",
		X"36",X"01",X"00",X"18",X"B4",X"21",X"BB",X"F0",X"35",X"28",X"10",X"2A",X"81",X"F0",X"ED",X"5B",
		X"85",X"F0",X"19",X"7C",X"DD",X"86",X"03",X"DD",X"77",X"03",X"C9",X"36",X"03",X"AF",X"DD",X"77",
		X"00",X"32",X"BE",X"F0",X"FD",X"2A",X"BF",X"F0",X"FD",X"36",X"02",X"A2",X"18",X"8B",X"21",X"BB",
		X"F0",X"35",X"C0",X"FD",X"2A",X"BF",X"F0",X"FD",X"36",X"02",X"75",X"AF",X"32",X"BA",X"F0",X"21",
		X"8E",X"F3",X"3E",X"10",X"96",X"30",X"01",X"AF",X"32",X"BB",X"F0",X"C9",X"3A",X"C2",X"F0",X"B7",
		X"C4",X"1D",X"3A",X"3A",X"C1",X"F0",X"B7",X"28",X"17",X"DD",X"21",X"D8",X"F8",X"21",X"5A",X"39",
		X"3D",X"47",X"CB",X"27",X"80",X"85",X"30",X"01",X"24",X"6F",X"E9",X"21",X"C1",X"F0",X"34",X"C9",
		X"3A",X"C3",X"F0",X"B7",X"C8",X"3D",X"32",X"C3",X"F0",X"C9",X"C3",X"60",X"39",X"C3",X"9C",X"39",
		X"21",X"C3",X"F0",X"35",X"28",X"23",X"FD",X"2A",X"CC",X"F0",X"3A",X"C4",X"F0",X"FD",X"86",X"05",
		X"DD",X"77",X"00",X"DD",X"7E",X"01",X"B7",X"3E",X"04",X"20",X"02",X"ED",X"44",X"21",X"C5",X"F0",
		X"86",X"77",X"FD",X"86",X"07",X"DD",X"77",X"03",X"C9",X"3E",X"04",X"77",X"32",X"C4",X"F0",X"CD",
		X"4B",X"39",X"FD",X"2A",X"C6",X"F0",X"DD",X"7E",X"01",X"FD",X"77",X"01",X"FD",X"2A",X"CC",X"F0",
		X"CD",X"73",X"39",X"FD",X"2A",X"C6",X"F0",X"21",X"C3",X"F0",X"35",X"28",X"14",X"86",X"C6",X"04",
		X"FD",X"77",X"03",X"3A",X"C4",X"F0",X"3D",X"32",X"C4",X"F0",X"DD",X"86",X"00",X"FD",X"77",X"00",
		X"C9",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"FD",X"36",X"02",
		X"A9",X"AF",X"DD",X"77",X"00",X"32",X"C1",X"F0",X"3A",X"C2",X"F0",X"B7",X"20",X"05",X"0E",X"2F",
		X"CD",X"4E",X"3D",X"3C",X"32",X"C2",X"F0",X"21",X"8E",X"F3",X"3E",X"10",X"96",X"30",X"01",X"AF",
		X"32",X"C3",X"F0",X"FD",X"7E",X"01",X"B7",X"C0",X"FD",X"2A",X"CC",X"F0",X"FD",X"7E",X"01",X"E6",
		X"0A",X"C0",X"FD",X"7E",X"05",X"FE",X"80",X"3E",X"02",X"38",X"02",X"ED",X"44",X"FD",X"77",X"04",
		X"FD",X"36",X"0C",X"04",X"FD",X"7E",X"01",X"F6",X"04",X"FD",X"77",X"01",X"C9",X"16",X"02",X"DD",
		X"21",X"60",X"F8",X"21",X"C8",X"F0",X"DD",X"7E",X"00",X"B7",X"CA",X"FA",X"3A",X"DD",X"7E",X"02",
		X"FE",X"6C",X"CA",X"FA",X"3A",X"7E",X"FE",X"FF",X"CA",X"C6",X"3A",X"B7",X"3A",X"82",X"F0",X"28",
		X"1C",X"C6",X"02",X"DD",X"86",X"03",X"30",X"1C",X"DD",X"36",X"00",X"00",X"3A",X"C2",X"F0",X"3D",
		X"32",X"C2",X"F0",X"B7",X"C2",X"FA",X"3A",X"0E",X"4C",X"CD",X"4E",X"3D",X"C9",X"D6",X"0D",X"DD",
		X"86",X"03",X"30",X"E4",X"DD",X"77",X"03",X"E5",X"DD",X"7E",X"03",X"DD",X"86",X"01",X"4F",X"06",
		X"00",X"FD",X"21",X"5B",X"F2",X"CD",X"B5",X"41",X"E1",X"DD",X"7E",X"00",X"C6",X"08",X"FD",X"BE",
		X"00",X"38",X"15",X"FD",X"BE",X"01",X"38",X"2A",X"47",X"FD",X"7E",X"02",X"B7",X"28",X"09",X"B8",
		X"30",X"06",X"FD",X"7E",X"03",X"B8",X"30",X"1A",X"DD",X"36",X"02",X"39",X"36",X"FF",X"23",X"36",
		X"04",X"0E",X"4C",X"3A",X"C2",X"F0",X"FE",X"02",X"DC",X"4E",X"3D",X"0E",X"15",X"CD",X"4E",X"3D",
		X"18",X"48",X"23",X"35",X"20",X"44",X"36",X"02",X"0E",X"A9",X"DD",X"7E",X"02",X"B9",X"20",X"01",
		X"0C",X"DD",X"71",X"02",X"18",X"34",X"E5",X"2A",X"81",X"F0",X"ED",X"4B",X"85",X"F0",X"09",X"7C",
		X"E1",X"DD",X"86",X"03",X"38",X"19",X"DD",X"77",X"03",X"23",X"35",X"20",X"1D",X"36",X"04",X"DD",
		X"7E",X"02",X"FE",X"39",X"20",X"04",X"3E",X"A2",X"18",X"0D",X"3C",X"FE",X"A7",X"38",X"08",X"0E",
		X"16",X"CD",X"4E",X"3D",X"C3",X"48",X"3A",X"DD",X"77",X"02",X"15",X"C8",X"DD",X"21",X"64",X"F8",
		X"21",X"CA",X"F0",X"C3",X"26",X"3A",X"3A",X"15",X"F0",X"B7",X"DD",X"7E",X"02",X"28",X"07",X"E6",
		X"80",X"20",X"08",X"C3",X"32",X"3F",X"E6",X"80",X"C2",X"32",X"3F",X"DD",X"7E",X"0A",X"B7",X"28",
		X"08",X"FE",X"10",X"30",X"04",X"DD",X"35",X"0A",X"C9",X"DD",X"36",X"07",X"E8",X"CD",X"F3",X"43",
		X"FD",X"21",X"5B",X"F2",X"FD",X"7E",X"00",X"B7",X"C8",X"DD",X"36",X"07",X"F8",X"DD",X"7E",X"02",
		X"E6",X"0F",X"28",X"04",X"FE",X"06",X"38",X"4E",X"47",X"DD",X"7E",X"09",X"FE",X"FF",X"20",X"4D",
		X"3A",X"06",X"F0",X"FE",X"01",X"20",X"0F",X"FD",X"7E",X"02",X"B7",X"28",X"0D",X"FD",X"77",X"00",
		X"FD",X"7E",X"03",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"DD",X"7E",X"01",X"E6",X"01",X"28",
		X"42",X"3A",X"06",X"F0",X"DD",X"77",X"09",X"78",X"B7",X"20",X"13",X"3A",X"06",X"F0",X"FE",X"02",
		X"30",X"0C",X"CB",X"42",X"28",X"08",X"FD",X"7E",X"01",X"D6",X"02",X"C3",X"B3",X"3C",X"FD",X"7E",
		X"00",X"D6",X"0E",X"C3",X"B3",X"3C",X"DD",X"7E",X"09",X"FE",X"FF",X"28",X"16",X"B7",X"28",X"0F",
		X"FD",X"7E",X"02",X"B7",X"28",X"0D",X"FD",X"77",X"00",X"FD",X"7E",X"03",X"FD",X"77",X"01",X"FD",
		X"36",X"02",X"00",X"1E",X"00",X"FD",X"21",X"8B",X"F2",X"7B",X"FE",X"06",X"CA",X"54",X"3C",X"FD",
		X"7E",X"00",X"DD",X"BE",X"00",X"CA",X"4B",X"3C",X"FD",X"7E",X"05",X"B7",X"28",X"7D",X"DD",X"7E",
		X"10",X"FD",X"96",X"10",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"47",X"DD",X"7E",X"08",X"B7",X"20",
		X"16",X"FD",X"B6",X"08",X"20",X"65",X"78",X"ED",X"44",X"FD",X"86",X"0E",X"FD",X"86",X"07",X"38",
		X"17",X"FE",X"F0",X"30",X"13",X"18",X"54",X"FD",X"7E",X"08",X"B7",X"20",X"0B",X"FD",X"7E",X"07",
		X"90",X"38",X"05",X"DD",X"BE",X"0E",X"30",X"43",X"DD",X"E5",X"DD",X"21",X"66",X"F2",X"DD",X"36",
		X"00",X"10",X"FD",X"7E",X"05",X"DD",X"77",X"01",X"C6",X"10",X"DD",X"77",X"02",X"DD",X"36",X"03",
		X"F0",X"DD",X"36",X"04",X"00",X"FD",X"E5",X"DD",X"E5",X"DD",X"21",X"5B",X"F2",X"FD",X"21",X"71",
		X"F2",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",X"23",X"FD",X"23",X"B7",X"20",X"F3",X"DD",X"E1",
		X"FD",X"21",X"71",X"F2",X"CD",X"DE",X"44",X"FD",X"E1",X"DD",X"E1",X"01",X"23",X"00",X"FD",X"09",
		X"1C",X"C3",X"B9",X"3B",X"FD",X"21",X"5B",X"F2",X"FD",X"7E",X"00",X"B7",X"C8",X"DD",X"7E",X"0A",
		X"B7",X"28",X"0E",X"47",X"CD",X"62",X"45",X"30",X"03",X"78",X"18",X"47",X"DD",X"36",X"0A",X"0F",
		X"C9",X"CD",X"E7",X"3C",X"47",X"FD",X"7E",X"02",X"B7",X"28",X"20",X"FD",X"7E",X"04",X"B7",X"28",
		X"0D",X"78",X"CB",X"47",X"28",X"08",X"FD",X"7E",X"05",X"FD",X"5E",X"04",X"18",X"13",X"78",X"CB",
		X"4F",X"28",X"08",X"FD",X"7E",X"03",X"FD",X"5E",X"02",X"18",X"06",X"FD",X"7E",X"01",X"FD",X"5E",
		X"00",X"93",X"D6",X"20",X"D8",X"28",X"09",X"4F",X"78",X"B9",X"38",X"04",X"CB",X"3F",X"18",X"F9",
		X"83",X"C6",X"08",X"DD",X"77",X"05",X"DD",X"7E",X"01",X"EE",X"10",X"DD",X"77",X"01",X"DD",X"7E",
		X"02",X"47",X"E6",X"10",X"C8",X"DD",X"7E",X"08",X"B7",X"28",X"04",X"DD",X"36",X"07",X"E8",X"78",
		X"E6",X"0F",X"C0",X"DD",X"36",X"0D",X"01",X"AF",X"32",X"4B",X"F0",X"32",X"4C",X"F0",X"DD",X"7E",
		X"01",X"E6",X"01",X"32",X"4A",X"F0",X"C9",X"3A",X"00",X"F4",X"07",X"30",X"02",X"EE",X"2B",X"C5",
		X"47",X"ED",X"5F",X"A8",X"C1",X"32",X"00",X"F4",X"C9",X"3A",X"8F",X"F3",X"D3",X"E0",X"FE",X"01",
		X"38",X"F7",X"AF",X"32",X"8F",X"F3",X"C9",X"06",X"10",X"DD",X"21",X"00",X"FA",X"11",X"02",X"00",
		X"7E",X"B7",X"28",X"03",X"1B",X"DD",X"23",X"23",X"7E",X"DD",X"77",X"00",X"DD",X"77",X"40",X"23",
		X"DD",X"19",X"10",X"E9",X"C9",X"21",X"91",X"F3",X"C3",X"2E",X"3D",X"21",X"2A",X"F4",X"2D",X"36",
		X"00",X"20",X"FB",X"25",X"7C",X"FE",X"F0",X"30",X"F5",X"C9",X"21",X"04",X"F8",X"06",X"7F",X"36",
		X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"36",X"00",X"23",X"10",X"F2",X"C9",X"F3",X"F5",
		X"3A",X"18",X"F4",X"B7",X"79",X"20",X"0F",X"FE",X"09",X"30",X"30",X"FE",X"02",X"20",X"0F",X"3E",
		X"01",X"32",X"18",X"F4",X"18",X"08",X"FE",X"01",X"20",X"04",X"AF",X"32",X"18",X"F4",X"3A",X"1D",
		X"F4",X"FE",X"0C",X"30",X"16",X"3C",X"32",X"1D",X"F4",X"E5",X"2A",X"1B",X"F4",X"CB",X"79",X"28",
		X"04",X"79",X"E6",X"7F",X"4F",X"71",X"23",X"22",X"1B",X"F4",X"E1",X"F1",X"FB",X"C9",X"F3",X"F5",
		X"E5",X"3A",X"18",X"F4",X"B7",X"28",X"18",X"3A",X"1D",X"F4",X"C6",X"03",X"FE",X"0C",X"30",X"0F",
		X"32",X"1D",X"F4",X"2A",X"1B",X"F4",X"71",X"23",X"72",X"23",X"73",X"23",X"22",X"1B",X"F4",X"E1",
		X"F1",X"FB",X"C9",X"C5",X"D5",X"FD",X"21",X"04",X"F8",X"11",X"04",X"00",X"06",X"14",X"3A",X"15",
		X"F0",X"B7",X"28",X"02",X"06",X"11",X"48",X"FD",X"7E",X"00",X"B7",X"28",X"0B",X"FD",X"19",X"10",
		X"F6",X"FD",X"21",X"04",X"F8",X"AF",X"18",X"09",X"3A",X"AD",X"F0",X"3C",X"32",X"AD",X"F0",X"79",
		X"90",X"D1",X"C1",X"C9",X"21",X"41",X"F1",X"85",X"30",X"01",X"24",X"6F",X"7E",X"C9",X"3A",X"28",
		X"F0",X"B7",X"C0",X"C5",X"FD",X"E5",X"E5",X"FD",X"E1",X"21",X"88",X"F3",X"06",X"06",X"7E",X"0E",
		X"00",X"FD",X"86",X"06",X"30",X"05",X"0C",X"C6",X"06",X"18",X"07",X"FE",X"0A",X"38",X"03",X"0C",
		X"D6",X"0A",X"77",X"2B",X"FD",X"2B",X"79",X"B7",X"28",X"01",X"34",X"10",X"E1",X"3A",X"8A",X"F2",
		X"B7",X"28",X"3B",X"21",X"88",X"F3",X"FD",X"21",X"82",X"F2",X"06",X"06",X"7E",X"FD",X"BE",X"00",
		X"38",X"2C",X"2B",X"FD",X"2B",X"10",X"F5",X"21",X"8A",X"F2",X"35",X"C4",X"62",X"3E",X"21",X"89",
		X"F3",X"7E",X"34",X"0E",X"0B",X"CD",X"4E",X"3D",X"FE",X"08",X"30",X"12",X"ED",X"44",X"21",X"70",
		X"E8",X"85",X"6F",X"06",X"01",X"3A",X"14",X"F0",X"B7",X"28",X"02",X"06",X"76",X"70",X"FD",X"E1",
		X"C1",X"C9",X"C5",X"FD",X"E5",X"FD",X"21",X"83",X"F2",X"21",X"82",X"F2",X"06",X"06",X"7E",X"0E",
		X"00",X"FD",X"86",X"06",X"30",X"05",X"0C",X"C6",X"06",X"18",X"07",X"FE",X"0A",X"38",X"03",X"0C",
		X"D6",X"0A",X"77",X"2B",X"FD",X"2B",X"79",X"B7",X"28",X"01",X"34",X"10",X"E1",X"FD",X"E1",X"C1",
		X"C9",X"E6",X"0F",X"28",X"56",X"FE",X"02",X"38",X"25",X"21",X"28",X"F0",X"3A",X"8E",X"F3",X"3C",
		X"CB",X"27",X"C6",X"08",X"86",X"77",X"3A",X"5E",X"F0",X"B7",X"28",X"18",X"AF",X"32",X"5E",X"F0",
		X"3A",X"5D",X"F0",X"B7",X"20",X"0E",X"3A",X"12",X"F0",X"EE",X"04",X"32",X"12",X"F0",X"21",X"52",
		X"B9",X"CD",X"EE",X"3D",X"3A",X"49",X"F0",X"B7",X"C0",X"21",X"45",X"F0",X"7E",X"B7",X"C0",X"3A",
		X"15",X"F0",X"B7",X"0E",X"01",X"20",X"02",X"0E",X"0A",X"7B",X"E6",X"03",X"CB",X"27",X"81",X"77",
		X"79",X"B3",X"CB",X"47",X"C0",X"21",X"42",X"F0",X"36",X"01",X"C9",X"21",X"59",X"B9",X"CD",X"EE",
		X"3D",X"3A",X"8E",X"F3",X"FE",X"02",X"D8",X"21",X"E7",X"F0",X"7E",X"B7",X"C0",X"36",X"80",X"C9",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"00",X"11",X"00",X"3F",X"F3",X"C5",X"3A",X"14",X"F0",X"FE",X"01",X"0E",
		X"1B",X"28",X"02",X"0E",X"00",X"1A",X"B7",X"28",X"06",X"81",X"77",X"13",X"2B",X"18",X"F6",X"C1",
		X"FB",X"C9",X"C5",X"E5",X"0E",X"00",X"DD",X"7E",X"18",X"B7",X"28",X"08",X"DD",X"71",X"18",X"67",
		X"DD",X"6E",X"17",X"71",X"DD",X"7E",X"13",X"B7",X"28",X"08",X"DD",X"71",X"13",X"67",X"DD",X"6E",
		X"12",X"71",X"DD",X"7E",X"15",X"B7",X"28",X"08",X"DD",X"71",X"15",X"67",X"DD",X"6E",X"14",X"71",
		X"DD",X"71",X"05",X"DD",X"71",X"01",X"21",X"32",X"F0",X"35",X"DD",X"7E",X"02",X"E6",X"0F",X"C2",
		X"7D",X"3F",X"32",X"49",X"F0",X"32",X"46",X"F0",X"CD",X"01",X"56",X"18",X"18",X"FE",X"06",X"38",
		X"14",X"AF",X"32",X"58",X"F0",X"32",X"60",X"F0",X"3A",X"33",X"F0",X"FE",X"03",X"20",X"06",X"3A",
		X"34",X"F0",X"32",X"33",X"F0",X"E1",X"C1",X"C9",X"C5",X"D5",X"FD",X"21",X"00",X"F9",X"11",X"04",
		X"00",X"06",X"30",X"3A",X"9E",X"F0",X"B7",X"28",X"02",X"06",X"2A",X"48",X"FD",X"7E",X"00",X"B7",
		X"28",X"1C",X"FD",X"19",X"10",X"F6",X"CD",X"E7",X"3C",X"E6",X"1F",X"47",X"CB",X"27",X"CB",X"27",
		X"11",X"00",X"F9",X"83",X"30",X"01",X"14",X"5F",X"D5",X"FD",X"E1",X"78",X"18",X"09",X"3A",X"D8",
		X"F0",X"3C",X"32",X"D8",X"F0",X"79",X"90",X"D1",X"C1",X"C9",X"21",X"0B",X"F1",X"85",X"30",X"01",
		X"24",X"6F",X"7E",X"C9",X"FD",X"21",X"5B",X"F2",X"C5",X"06",X"00",X"0E",X"00",X"CD",X"B5",X"41",
		X"FD",X"7E",X"00",X"B7",X"28",X"5E",X"CD",X"E7",X"3C",X"47",X"FD",X"7E",X"02",X"B7",X"28",X"0C",
		X"CB",X"48",X"28",X"08",X"FD",X"7E",X"03",X"FD",X"5E",X"02",X"18",X"06",X"FD",X"7E",X"01",X"FD",
		X"5E",X"00",X"93",X"D6",X"28",X"38",X"3D",X"28",X"09",X"4F",X"78",X"B9",X"38",X"04",X"CB",X"3F",
		X"18",X"F9",X"83",X"C6",X"04",X"4F",X"CD",X"B3",X"3D",X"CD",X"E4",X"3D",X"36",X"01",X"FD",X"71",
		X"00",X"FD",X"36",X"03",X"00",X"FD",X"36",X"02",X"1E",X"CD",X"B3",X"3D",X"CD",X"E4",X"3D",X"36",
		X"02",X"CD",X"E7",X"3C",X"E6",X"07",X"C6",X"03",X"81",X"FD",X"77",X"00",X"FD",X"36",X"03",X"00",
		X"FD",X"36",X"02",X"1F",X"C1",X"C9",X"3A",X"01",X"F0",X"FE",X"B0",X"D0",X"DD",X"7E",X"01",X"E6",
		X"40",X"C0",X"DD",X"7E",X"02",X"E6",X"60",X"C8",X"C5",X"47",X"CD",X"CD",X"40",X"38",X"5C",X"21",
		X"51",X"F0",X"7E",X"B7",X"20",X"05",X"0E",X"31",X"CD",X"4E",X"3D",X"34",X"DD",X"7E",X"01",X"F6",
		X"40",X"DD",X"77",X"01",X"CB",X"68",X"28",X"26",X"FD",X"E5",X"D1",X"DD",X"73",X"12",X"DD",X"72",
		X"13",X"FD",X"36",X"00",X"01",X"FD",X"36",X"02",X"0D",X"FD",X"36",X"01",X"20",X"DD",X"7E",X"02",
		X"EE",X"20",X"DD",X"77",X"02",X"CB",X"70",X"28",X"22",X"CD",X"CD",X"40",X"38",X"1D",X"FD",X"E5",
		X"D1",X"DD",X"73",X"14",X"DD",X"72",X"15",X"FD",X"36",X"00",X"01",X"FD",X"36",X"02",X"0D",X"FD",
		X"36",X"01",X"00",X"DD",X"7E",X"02",X"EE",X"40",X"DD",X"77",X"02",X"C1",X"C9",X"0E",X"06",X"FD",
		X"21",X"90",X"F8",X"11",X"04",X"00",X"FD",X"7E",X"00",X"B7",X"C8",X"FD",X"19",X"0D",X"20",X"F6",
		X"37",X"C9",X"3A",X"BA",X"F0",X"21",X"BB",X"F0",X"B6",X"C0",X"DD",X"7E",X"07",X"FE",X"08",X"D8",
		X"DD",X"7E",X"18",X"B7",X"C8",X"67",X"DD",X"6E",X"17",X"22",X"BD",X"F0",X"AF",X"DD",X"77",X"18",
		X"3C",X"32",X"BA",X"F0",X"DD",X"7E",X"10",X"C6",X"04",X"32",X"BC",X"F0",X"21",X"BB",X"F0",X"36",
		X"06",X"C9",X"3A",X"C1",X"F0",X"21",X"C3",X"F0",X"B6",X"C0",X"DD",X"7E",X"07",X"FE",X"08",X"D8",
		X"FE",X"E4",X"D0",X"DD",X"7E",X"18",X"B7",X"C8",X"16",X"00",X"FD",X"21",X"60",X"F8",X"FD",X"7E",
		X"00",X"B7",X"28",X"0C",X"14",X"FD",X"21",X"64",X"F8",X"FD",X"7E",X"00",X"B7",X"28",X"01",X"C9",
		X"FD",X"22",X"C6",X"F0",X"FD",X"36",X"00",X"01",X"FD",X"36",X"02",X"6C",X"DD",X"22",X"CC",X"F0",
		X"C5",X"06",X"00",X"3A",X"01",X"F0",X"DD",X"BE",X"07",X"38",X"02",X"06",X"10",X"21",X"C8",X"F0",
		X"7A",X"CB",X"27",X"85",X"30",X"01",X"24",X"6F",X"70",X"23",X"36",X"04",X"7B",X"B7",X"3E",X"06",
		X"20",X"02",X"3E",X"F9",X"32",X"C4",X"F0",X"FD",X"21",X"D8",X"F8",X"DD",X"86",X"05",X"FD",X"77",
		X"00",X"3E",X"09",X"32",X"C5",X"F0",X"DD",X"86",X"07",X"FD",X"77",X"03",X"FD",X"70",X"01",X"FD",
		X"36",X"02",X"A8",X"3E",X"01",X"32",X"C1",X"F0",X"21",X"C3",X"F0",X"36",X"03",X"0E",X"4D",X"CD",
		X"4E",X"3D",X"3A",X"8E",X"F3",X"CB",X"27",X"CB",X"27",X"47",X"3E",X"40",X"90",X"30",X"01",X"AF",
		X"DD",X"77",X"1C",X"C1",X"C9",X"DD",X"E5",X"CD",X"5A",X"4B",X"DD",X"7E",X"00",X"32",X"54",X"F0",
		X"E6",X"0F",X"6F",X"CB",X"27",X"85",X"21",X"D2",X"41",X"85",X"30",X"01",X"24",X"6F",X"DD",X"7E",
		X"01",X"E9",X"C3",X"02",X"42",X"C3",X"0E",X"42",X"C3",X"41",X"42",X"C3",X"53",X"42",X"C3",X"62",
		X"42",X"C3",X"80",X"42",X"C3",X"A0",X"42",X"C3",X"BE",X"42",X"C3",X"DC",X"42",X"C3",X"0C",X"43",
		X"C3",X"3E",X"43",X"C3",X"70",X"43",X"C3",X"8C",X"43",X"C3",X"AC",X"43",X"C3",X"CE",X"43",X"C3",
		X"E4",X"43",X"F5",X"3A",X"15",X"F0",X"B7",X"C2",X"45",X"43",X"F1",X"C3",X"53",X"42",X"3A",X"15",
		X"F0",X"B7",X"20",X"18",X"DD",X"7E",X"01",X"C6",X"10",X"DD",X"86",X"02",X"FD",X"77",X"00",X"DD",
		X"86",X"03",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"C3",X"F0",X"43",X"DD",X"7E",X"01",X"C6",
		X"10",X"FD",X"77",X"00",X"DD",X"86",X"02",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"C3",X"F0",
		X"43",X"C6",X"10",X"FD",X"77",X"00",X"DD",X"86",X"02",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",
		X"C3",X"F0",X"43",X"FD",X"36",X"00",X"92",X"FD",X"36",X"01",X"E2",X"FD",X"36",X"02",X"00",X"C3",
		X"F0",X"43",X"C6",X"10",X"FD",X"77",X"00",X"DD",X"86",X"02",X"FD",X"77",X"01",X"DD",X"86",X"03",
		X"FD",X"77",X"02",X"DD",X"86",X"02",X"FD",X"77",X"03",X"FD",X"36",X"04",X"00",X"C3",X"F0",X"43",
		X"C6",X"10",X"FD",X"77",X"00",X"DD",X"86",X"02",X"FD",X"77",X"01",X"C6",X"20",X"DD",X"86",X"03",
		X"FD",X"77",X"02",X"DD",X"86",X"02",X"FD",X"77",X"03",X"FD",X"36",X"04",X"00",X"C3",X"F0",X"43",
		X"C6",X"10",X"FD",X"77",X"01",X"C6",X"20",X"DD",X"86",X"02",X"FD",X"77",X"02",X"DD",X"86",X"03",
		X"FD",X"77",X"03",X"FD",X"36",X"00",X"01",X"FD",X"36",X"04",X"00",X"C3",X"F0",X"43",X"C6",X"10",
		X"FD",X"77",X"00",X"DD",X"86",X"02",X"FD",X"77",X"01",X"C6",X"20",X"DD",X"86",X"03",X"FD",X"77",
		X"02",X"FD",X"36",X"03",X"FF",X"FD",X"36",X"04",X"00",X"C3",X"F0",X"43",X"F5",X"3A",X"15",X"F0",
		X"B7",X"28",X"13",X"F1",X"C6",X"10",X"FD",X"77",X"00",X"DD",X"86",X"02",X"FD",X"77",X"01",X"FD",
		X"36",X"02",X"00",X"C3",X"F0",X"43",X"F1",X"DD",X"86",X"02",X"C6",X"20",X"FD",X"77",X"00",X"DD",
		X"86",X"03",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"C3",X"F0",X"43",X"F5",X"3A",X"15",X"F0",
		X"B7",X"28",X"15",X"F1",X"C6",X"08",X"FD",X"77",X"00",X"DD",X"86",X"02",X"C6",X"10",X"FD",X"77",
		X"01",X"FD",X"36",X"02",X"00",X"C3",X"F0",X"43",X"F1",X"DD",X"86",X"02",X"C6",X"30",X"FD",X"77",
		X"00",X"DD",X"86",X"03",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"C3",X"F0",X"43",X"F5",X"3A",
		X"15",X"F0",X"B7",X"28",X"15",X"F1",X"C6",X"08",X"FD",X"77",X"00",X"DD",X"86",X"02",X"C6",X"10",
		X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"C3",X"F0",X"43",X"F1",X"DD",X"86",X"02",X"C6",X"50",
		X"FD",X"77",X"00",X"DD",X"86",X"03",X"FD",X"77",X"01",X"FD",X"36",X"02",X"00",X"C3",X"F0",X"43",
		X"C6",X"10",X"FD",X"77",X"00",X"DD",X"86",X"02",X"FD",X"77",X"01",X"C6",X"10",X"FD",X"77",X"02",
		X"DD",X"86",X"03",X"FD",X"77",X"03",X"FD",X"36",X"04",X"00",X"18",X"64",X"C6",X"08",X"FD",X"77",
		X"00",X"DD",X"86",X"02",X"C6",X"10",X"FD",X"77",X"01",X"C6",X"10",X"FD",X"77",X"02",X"DD",X"86",
		X"03",X"C6",X"10",X"FD",X"77",X"03",X"FD",X"36",X"04",X"00",X"18",X"44",X"C6",X"08",X"FD",X"77",
		X"00",X"DD",X"86",X"02",X"C6",X"10",X"FD",X"77",X"01",X"C6",X"20",X"C6",X"10",X"FD",X"77",X"02",
		X"DD",X"86",X"03",X"C6",X"10",X"FD",X"77",X"03",X"FD",X"36",X"04",X"00",X"18",X"22",X"B7",X"20",
		X"05",X"FD",X"77",X"00",X"18",X"1A",X"FD",X"36",X"00",X"3C",X"FD",X"36",X"01",X"7C",X"FD",X"36",
		X"02",X"00",X"18",X"0C",X"F5",X"3A",X"15",X"F0",X"B7",X"C2",X"45",X"43",X"F1",X"C3",X"53",X"42",
		X"DD",X"E1",X"C9",X"DD",X"E5",X"DD",X"46",X"08",X"DD",X"4E",X"07",X"FD",X"21",X"66",X"F2",X"CD",
		X"B5",X"41",X"3A",X"54",X"F0",X"32",X"55",X"F0",X"79",X"DD",X"86",X"0E",X"30",X"01",X"04",X"4F",
		X"FD",X"21",X"71",X"F2",X"CD",X"B5",X"41",X"3A",X"54",X"F0",X"E6",X"F0",X"21",X"55",X"F0",X"B6",
		X"77",X"DD",X"21",X"66",X"F2",X"CD",X"DE",X"44",X"DD",X"E1",X"DD",X"7E",X"08",X"B7",X"C0",X"3A",
		X"AD",X"F0",X"B7",X"C8",X"CB",X"7F",X"C0",X"4F",X"D5",X"11",X"04",X"00",X"FD",X"21",X"04",X"F8",
		X"06",X"00",X"FD",X"7E",X"00",X"B7",X"CA",X"CC",X"44",X"FE",X"E8",X"30",X"7C",X"78",X"CD",X"E4",
		X"3D",X"E6",X"0F",X"FE",X"03",X"38",X"72",X"6F",X"DD",X"7E",X"10",X"ED",X"44",X"CB",X"27",X"CB",
		X"27",X"CB",X"27",X"C6",X"28",X"FD",X"86",X"03",X"38",X"5F",X"DD",X"BE",X"07",X"38",X"5A",X"DD",
		X"7E",X"0E",X"CB",X"3F",X"DD",X"86",X"07",X"FD",X"BE",X"03",X"38",X"4D",X"DD",X"E5",X"FD",X"E5",
		X"DD",X"21",X"66",X"F2",X"7D",X"CB",X"27",X"CB",X"27",X"21",X"4D",X"BB",X"85",X"30",X"01",X"24",
		X"6F",X"DD",X"36",X"00",X"08",X"FD",X"7E",X"00",X"86",X"D6",X"04",X"DD",X"77",X"01",X"C6",X"08",
		X"23",X"86",X"DD",X"77",X"02",X"DD",X"36",X"03",X"FF",X"DD",X"36",X"04",X"00",X"FD",X"21",X"71",
		X"F2",X"21",X"5B",X"F2",X"7E",X"FD",X"77",X"00",X"23",X"FD",X"23",X"B7",X"20",X"F6",X"FD",X"21",
		X"71",X"F2",X"CD",X"DE",X"44",X"FD",X"E1",X"DD",X"E1",X"0D",X"28",X"10",X"FD",X"19",X"04",X"78",
		X"FE",X"14",X"C2",X"42",X"44",X"3A",X"AD",X"F0",X"0D",X"32",X"AD",X"F0",X"D1",X"C9",X"D5",X"21",
		X"5B",X"F2",X"01",X"02",X"00",X"DD",X"7E",X"00",X"B7",X"28",X"73",X"FD",X"7E",X"00",X"B7",X"28",
		X"6D",X"DD",X"7E",X"00",X"FD",X"BE",X"01",X"30",X"5D",X"FD",X"7E",X"00",X"DD",X"BE",X"01",X"30",
		X"59",X"DD",X"BE",X"00",X"30",X"03",X"DD",X"7E",X"00",X"77",X"FD",X"7E",X"01",X"DD",X"BE",X"01",
		X"30",X"1D",X"5F",X"96",X"D6",X"16",X"38",X"03",X"23",X"73",X"23",X"FD",X"09",X"FD",X"7E",X"00",
		X"DD",X"BE",X"01",X"38",X"C0",X"DD",X"7E",X"02",X"B7",X"28",X"BA",X"DD",X"09",X"18",X"B6",X"DD",
		X"7E",X"01",X"5F",X"FE",X"FF",X"28",X"0C",X"96",X"38",X"0C",X"D6",X"16",X"30",X"05",X"7E",X"FE",
		X"01",X"20",X"03",X"23",X"73",X"23",X"DD",X"09",X"DD",X"7E",X"00",X"FD",X"BE",X"01",X"38",X"95",
		X"FD",X"7E",X"02",X"B7",X"28",X"8F",X"FD",X"09",X"18",X"8B",X"DD",X"09",X"18",X"87",X"36",X"00",
		X"D1",X"C9",X"0E",X"00",X"FD",X"7E",X"00",X"B7",X"C8",X"90",X"D0",X"78",X"C6",X"10",X"30",X"02",
		X"3E",X"FF",X"FD",X"96",X"01",X"D8",X"3C",X"4F",X"FD",X"7E",X"02",X"B7",X"C8",X"90",X"38",X"06",
		X"B9",X"D0",X"0E",X"00",X"3F",X"C9",X"78",X"C6",X"10",X"30",X"02",X"3E",X"FF",X"FD",X"96",X"03",
		X"0E",X"01",X"D8",X"3C",X"4F",X"FD",X"7E",X"04",X"B7",X"C8",X"90",X"38",X"06",X"B9",X"D0",X"0E",
		X"00",X"3F",X"C9",X"78",X"C6",X"10",X"FD",X"96",X"05",X"4F",X"C9",X"3A",X"32",X"F0",X"B7",X"C8",
		X"FD",X"E5",X"C5",X"D5",X"E5",X"1E",X"00",X"FD",X"21",X"8B",X"F2",X"7B",X"FE",X"06",X"28",X"7B",
		X"FD",X"7E",X"05",X"B7",X"28",X"6D",X"FD",X"7E",X"08",X"B7",X"20",X"08",X"3A",X"01",X"F0",X"FD",
		X"BE",X"07",X"38",X"5F",X"FD",X"7E",X"07",X"FD",X"86",X"0E",X"DD",X"BE",X"03",X"38",X"54",X"DD",
		X"7E",X"03",X"C6",X"10",X"FD",X"BE",X"07",X"38",X"4A",X"DD",X"7E",X"00",X"C6",X"0A",X"FD",X"BE",
		X"05",X"38",X"40",X"FD",X"7E",X"05",X"C6",X"10",X"D6",X"06",X"DD",X"BE",X"00",X"38",X"34",X"FD",
		X"7E",X"06",X"FE",X"7C",X"20",X"07",X"0E",X"37",X"CD",X"4E",X"3D",X"18",X"20",X"FD",X"7E",X"01",
		X"47",X"E6",X"0A",X"20",X"18",X"78",X"F6",X"0A",X"FD",X"77",X"01",X"FD",X"36",X"16",X"00",X"FD",
		X"36",X"20",X"20",X"FD",X"7E",X"02",X"CD",X"91",X"3E",X"FD",X"36",X"0C",X"01",X"E1",X"36",X"00",
		X"37",X"18",X"09",X"01",X"23",X"00",X"FD",X"09",X"1C",X"18",X"80",X"E1",X"D1",X"C1",X"FD",X"E1",
		X"C9",X"3A",X"01",X"F4",X"B7",X"C0",X"21",X"5B",X"F1",X"3A",X"89",X"F0",X"85",X"30",X"01",X"24",
		X"6F",X"3A",X"8A",X"F0",X"B7",X"28",X"10",X"3D",X"32",X"8A",X"F0",X"DD",X"7E",X"FC",X"77",X"23",
		X"DD",X"7E",X"FD",X"77",X"C3",X"F3",X"46",X"3A",X"8B",X"F0",X"B7",X"28",X"19",X"3D",X"32",X"8B",
		X"F0",X"FD",X"2A",X"8C",X"F0",X"11",X"04",X"00",X"FD",X"19",X"FD",X"22",X"8C",X"F0",X"FD",X"E5",
		X"D1",X"73",X"23",X"72",X"18",X"6D",X"DD",X"7E",X"01",X"B7",X"20",X"26",X"DD",X"B6",X"00",X"20",
		X"0F",X"CD",X"6C",X"49",X"CD",X"DF",X"49",X"DD",X"2A",X"93",X"F0",X"DD",X"7E",X"01",X"18",X"12",
		X"DD",X"7E",X"00",X"3D",X"32",X"8A",X"F0",X"DD",X"7E",X"FE",X"77",X"23",X"DD",X"7E",X"FF",X"77",
		X"18",X"3D",X"FE",X"01",X"20",X"1D",X"DD",X"7E",X"00",X"3D",X"32",X"8B",X"F0",X"FD",X"21",X"8C",
		X"F0",X"DD",X"7E",X"FE",X"FD",X"77",X"00",X"DD",X"7E",X"FF",X"FD",X"77",X"01",X"DD",X"23",X"DD",
		X"23",X"18",X"9E",X"DD",X"5E",X"00",X"73",X"23",X"DD",X"56",X"01",X"72",X"1A",X"B7",X"20",X"0F",
		X"3A",X"9E",X"F0",X"B7",X"20",X"09",X"3C",X"32",X"9E",X"F0",X"21",X"9D",X"F0",X"36",X"6F",X"DD",
		X"23",X"DD",X"23",X"3A",X"89",X"F0",X"C6",X"02",X"32",X"89",X"F0",X"3A",X"9E",X"F0",X"B7",X"CA",
		X"15",X"48",X"FE",X"03",X"38",X"74",X"20",X"41",X"3A",X"15",X"F0",X"B7",X"28",X"33",X"3A",X"00",
		X"F0",X"FE",X"80",X"38",X"2C",X"CD",X"B3",X"3D",X"CD",X"E4",X"3D",X"36",X"06",X"FD",X"22",X"B4",
		X"F0",X"FD",X"36",X"00",X"C1",X"FD",X"36",X"01",X"00",X"CD",X"E7",X"3C",X"E6",X"03",X"21",X"68",
		X"49",X"85",X"30",X"01",X"24",X"6F",X"7E",X"FD",X"77",X"02",X"FD",X"36",X"03",X"06",X"C3",X"11",
		X"48",X"3E",X"05",X"32",X"9E",X"F0",X"C3",X"15",X"48",X"FE",X"04",X"C2",X"15",X"48",X"FD",X"2A",
		X"B4",X"F0",X"FD",X"7E",X"03",X"D6",X"10",X"30",X"01",X"AF",X"F5",X"CD",X"B3",X"3D",X"CD",X"E4",
		X"3D",X"F1",X"36",X"06",X"FD",X"22",X"B6",X"F0",X"FD",X"36",X"00",X"C1",X"FD",X"36",X"01",X"00",
		X"FD",X"36",X"02",X"29",X"FD",X"77",X"03",X"C3",X"11",X"48",X"3A",X"9D",X"F0",X"3D",X"32",X"9D",
		X"F0",X"FE",X"02",X"D2",X"15",X"48",X"3A",X"15",X"F0",X"B7",X"3E",X"22",X"28",X"02",X"C6",X"8F",
		X"4F",X"C6",X"10",X"67",X"C6",X"10",X"6F",X"11",X"04",X"00",X"FD",X"21",X"A8",X"F9",X"3A",X"9D",
		X"F0",X"B7",X"20",X"3C",X"FD",X"7E",X"03",X"D6",X"10",X"30",X"01",X"AF",X"FD",X"21",X"B4",X"F9",
		X"FD",X"71",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"7E",X"FD",X"77",X"03",X"FD",X"19",
		X"FD",X"74",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"7F",X"FD",X"77",X"03",X"FD",X"19",
		X"FD",X"75",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"80",X"FD",X"77",X"03",X"18",X"31",
		X"FD",X"71",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"81",X"FD",X"36",X"03",X"02",X"FD",
		X"19",X"FD",X"74",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"82",X"FD",X"36",X"03",X"02",
		X"FD",X"19",X"FD",X"75",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"83",X"FD",X"36",X"03",
		X"02",X"21",X"9E",X"F0",X"34",X"3A",X"88",X"F0",X"EE",X"01",X"32",X"88",X"F0",X"C8",X"3A",X"7A",
		X"F3",X"FE",X"02",X"28",X"58",X"3A",X"09",X"F0",X"B7",X"20",X"3A",X"3A",X"06",X"F0",X"FE",X"02",
		X"28",X"33",X"3A",X"03",X"F0",X"E6",X"40",X"20",X"3A",X"3A",X"15",X"F0",X"B7",X"28",X"13",X"21",
		X"4B",X"B9",X"CD",X"EE",X"3D",X"3A",X"C2",X"F0",X"B7",X"20",X"28",X"0E",X"4C",X"CD",X"4E",X"3D",
		X"18",X"21",X"21",X"44",X"B9",X"CD",X"EE",X"3D",X"3A",X"51",X"F0",X"B7",X"20",X"15",X"0E",X"32",
		X"CD",X"4E",X"3D",X"18",X"0E",X"0E",X"1D",X"3A",X"56",X"F0",X"E6",X"80",X"28",X"02",X"0E",X"0F",
		X"CD",X"4E",X"3D",X"3A",X"28",X"F0",X"B7",X"28",X"04",X"3D",X"32",X"28",X"F0",X"21",X"A9",X"F0",
		X"7E",X"B7",X"28",X"6D",X"23",X"35",X"20",X"69",X"2B",X"36",X"00",X"21",X"AB",X"F0",X"36",X"01",
		X"2A",X"3E",X"F0",X"22",X"3C",X"F0",X"3A",X"15",X"F0",X"B7",X"20",X"1D",X"21",X"57",X"F0",X"36",
		X"04",X"3E",X"01",X"32",X"5B",X"F0",X"32",X"5E",X"F0",X"32",X"5D",X"F0",X"3E",X"04",X"32",X"5C",
		X"F0",X"3A",X"12",X"F0",X"F6",X"04",X"32",X"12",X"F0",X"3A",X"8E",X"F3",X"FE",X"07",X"30",X"24",
		X"3C",X"32",X"8E",X"F3",X"2A",X"30",X"F0",X"85",X"30",X"01",X"24",X"6F",X"7E",X"32",X"33",X"F0",
		X"3A",X"47",X"F0",X"CB",X"3F",X"32",X"47",X"F0",X"3A",X"40",X"F0",X"B7",X"28",X"13",X"3D",X"32",
		X"40",X"F0",X"18",X"0D",X"21",X"33",X"F0",X"36",X"06",X"FE",X"0C",X"30",X"04",X"3C",X"32",X"8E",
		X"F3",X"FD",X"21",X"61",X"F0",X"ED",X"5B",X"7A",X"F0",X"FD",X"19",X"FD",X"35",X"02",X"20",X"1A",
		X"FD",X"7E",X"01",X"21",X"33",X"F0",X"BE",X"38",X"01",X"7E",X"32",X"35",X"F0",X"7B",X"C6",X"03",
		X"FE",X"18",X"20",X"01",X"AF",X"5F",X"ED",X"53",X"7A",X"F0",X"0E",X"0F",X"FD",X"21",X"F2",X"DF",
		X"3A",X"16",X"F0",X"B7",X"28",X"05",X"11",X"00",X"04",X"FD",X"19",X"ED",X"5B",X"97",X"F0",X"FD",
		X"19",X"2A",X"95",X"F0",X"C5",X"7E",X"FE",X"44",X"28",X"04",X"FE",X"EF",X"20",X"0D",X"E6",X"BF",
		X"23",X"46",X"05",X"FD",X"77",X"00",X"FD",X"23",X"0D",X"10",X"F8",X"FD",X"77",X"00",X"23",X"FD",
		X"23",X"0D",X"20",X"E1",X"C1",X"22",X"95",X"F0",X"7B",X"D6",X"10",X"5F",X"30",X"05",X"7A",X"3D",
		X"E6",X"03",X"57",X"ED",X"53",X"97",X"F0",X"C9",X"6A",X"6B",X"69",X"6A",X"F5",X"3A",X"9F",X"F0",
		X"B7",X"28",X"24",X"3D",X"32",X"9F",X"F0",X"20",X"1E",X"C5",X"E5",X"21",X"A0",X"F0",X"36",X"01",
		X"0E",X"02",X"21",X"93",X"E9",X"06",X"0A",X"77",X"2B",X"10",X"FC",X"0D",X"28",X"07",X"21",X"15",
		X"EA",X"06",X"0E",X"18",X"F2",X"E1",X"C1",X"3A",X"E5",X"F0",X"B7",X"28",X"26",X"3A",X"E8",X"F0",
		X"B7",X"20",X"20",X"3A",X"E7",X"F0",X"B7",X"20",X"1A",X"CD",X"E7",X"3C",X"E5",X"21",X"E6",X"F0",
		X"BE",X"30",X"09",X"36",X"00",X"21",X"E7",X"F0",X"36",X"04",X"18",X"06",X"7E",X"C6",X"01",X"38",
		X"01",X"77",X"E1",X"F1",X"C9",X"42",X"52",X"49",X"44",X"47",X"45",X"20",X"4F",X"55",X"54",X"00",
		X"44",X"45",X"54",X"4F",X"55",X"52",X"20",X"4F",X"4E",X"20",X"4C",X"45",X"46",X"54",X"00",X"E5",
		X"C5",X"FD",X"E5",X"2A",X"99",X"F0",X"3A",X"8F",X"F0",X"B7",X"28",X"09",X"3D",X"32",X"8F",X"F0",
		X"3A",X"8E",X"F0",X"18",X"07",X"3A",X"90",X"F0",X"3C",X"32",X"90",X"F0",X"C6",X"02",X"CB",X"27",
		X"85",X"30",X"01",X"24",X"6F",X"E5",X"DD",X"E1",X"DD",X"7E",X"01",X"FE",X"01",X"D2",X"CC",X"4A",
		X"DD",X"B6",X"00",X"C2",X"BC",X"4A",X"21",X"99",X"F0",X"3A",X"15",X"F0",X"B7",X"20",X"17",X"3A",
		X"03",X"F0",X"E6",X"10",X"28",X"09",X"FD",X"2A",X"5F",X"F0",X"FD",X"7E",X"05",X"18",X"03",X"3A",
		X"00",X"F0",X"FE",X"80",X"30",X"0B",X"DD",X"7E",X"02",X"77",X"DD",X"7E",X"03",X"23",X"77",X"18",
		X"09",X"DD",X"7E",X"04",X"77",X"DD",X"7E",X"05",X"23",X"77",X"21",X"90",X"F0",X"36",X"00",X"DD",
		X"2A",X"99",X"F0",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"3A",X"15",X"F0",X"B7",X"20",X"19",X"3A",
		X"14",X"F0",X"B7",X"20",X"13",X"3A",X"8E",X"F3",X"FE",X"03",X"38",X"0C",X"57",X"CD",X"E7",X"3C",
		X"E6",X"0F",X"BA",X"30",X"03",X"21",X"83",X"C9",X"22",X"A7",X"F0",X"11",X"83",X"C9",X"7A",X"BC",
		X"20",X"1F",X"7B",X"BD",X"20",X"1B",X"21",X"8F",X"E9",X"11",X"27",X"B9",X"CD",X"18",X"3F",X"21",
		X"D0",X"E9",X"11",X"2B",X"B9",X"CD",X"18",X"3F",X"21",X"10",X"EA",X"11",X"31",X"B9",X"CD",X"18",
		X"3F",X"21",X"A9",X"F0",X"36",X"01",X"23",X"36",X"4E",X"DD",X"23",X"DD",X"23",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"22",X"3E",X"F0",X"DD",X"23",X"DD",X"23",X"18",X"3D",X"DD",X"7E",X"00",X"32",
		X"8F",X"F0",X"3A",X"90",X"F0",X"3D",X"32",X"8E",X"F0",X"C3",X"E3",X"49",X"20",X"2B",X"CD",X"E7",
		X"3C",X"E6",X"07",X"3C",X"21",X"8E",X"F3",X"96",X"21",X"6B",X"C0",X"30",X"22",X"21",X"93",X"E9",
		X"11",X"C5",X"49",X"CD",X"18",X"3F",X"21",X"15",X"EA",X"11",X"D0",X"49",X"CD",X"18",X"3F",X"21",
		X"9F",X"F0",X"36",X"04",X"21",X"A1",X"C3",X"18",X"06",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"5E",
		X"23",X"56",X"ED",X"53",X"95",X"F0",X"23",X"7E",X"01",X"03",X"00",X"ED",X"5B",X"7A",X"F0",X"FD",
		X"21",X"61",X"F0",X"FD",X"19",X"ED",X"5B",X"7C",X"F0",X"DD",X"21",X"61",X"F0",X"DD",X"19",X"DD",
		X"77",X"01",X"23",X"23",X"22",X"93",X"F0",X"2E",X"40",X"FD",X"7E",X"00",X"DD",X"BE",X"00",X"28",
		X"14",X"7D",X"FD",X"96",X"02",X"6F",X"FD",X"09",X"FD",X"7E",X"00",X"FE",X"08",X"20",X"EA",X"FD",
		X"21",X"61",X"F0",X"18",X"E4",X"DD",X"75",X"02",X"7B",X"C6",X"03",X"FE",X"18",X"20",X"01",X"AF",
		X"5F",X"ED",X"53",X"7C",X"F0",X"FD",X"E1",X"C1",X"E1",X"C9",X"FD",X"E5",X"C5",X"3A",X"15",X"F0",
		X"B7",X"28",X"07",X"79",X"D6",X"30",X"30",X"01",X"05",X"4F",X"FD",X"21",X"5B",X"F1",X"78",X"ED",
		X"44",X"47",X"79",X"ED",X"44",X"20",X"01",X"04",X"21",X"87",X"F0",X"86",X"F5",X"E6",X"F0",X"4F",
		X"F1",X"79",X"1F",X"1F",X"1F",X"4F",X"78",X"0F",X"0F",X"0F",X"30",X"01",X"79",X"A9",X"21",X"89",
		X"F0",X"86",X"C6",X"02",X"06",X"00",X"4F",X"FD",X"09",X"FD",X"6E",X"00",X"FD",X"66",X"01",X"E5",
		X"DD",X"E1",X"C1",X"FD",X"E1",X"C9",X"3A",X"38",X"F0",X"B7",X"28",X"04",X"3D",X"32",X"38",X"F0",
		X"16",X"00",X"DD",X"21",X"8B",X"F2",X"7A",X"FE",X"06",X"28",X"60",X"DD",X"7E",X"01",X"E6",X"80",
		X"28",X"05",X"CD",X"9C",X"0E",X"18",X"4C",X"DD",X"7E",X"01",X"B7",X"20",X"46",X"3A",X"32",X"F0",
		X"21",X"35",X"F0",X"BE",X"38",X"20",X"7E",X"B7",X"28",X"39",X"3A",X"06",X"F0",X"FE",X"02",X"30",
		X"32",X"3A",X"60",X"F0",X"B7",X"20",X"2C",X"3A",X"57",X"F0",X"FE",X"01",X"38",X"25",X"28",X"06",
		X"3D",X"32",X"57",X"F0",X"18",X"1D",X"3A",X"38",X"F0",X"B7",X"20",X"17",X"CD",X"E7",X"3C",X"E6",
		X"07",X"21",X"39",X"F0",X"86",X"2A",X"81",X"F0",X"CB",X"3C",X"CB",X"3C",X"94",X"32",X"38",X"F0",
		X"CD",X"76",X"0C",X"01",X"23",X"00",X"DD",X"09",X"14",X"18",X"9B",X"16",X"00",X"DD",X"21",X"8B",
		X"F2",X"7A",X"FE",X"06",X"C8",X"DD",X"7E",X"01",X"47",X"E6",X"10",X"28",X"05",X"CD",X"06",X"3B",
		X"18",X"06",X"78",X"E6",X"20",X"C4",X"23",X"14",X"01",X"23",X"00",X"DD",X"09",X"14",X"18",X"E1",
		X"DD",X"21",X"FF",X"F0",X"DD",X"7E",X"00",X"47",X"FE",X"01",X"DA",X"F0",X"51",X"28",X"7D",X"FE",
		X"02",X"28",X"69",X"FE",X"06",X"30",X"65",X"3A",X"E8",X"F0",X"B7",X"28",X"54",X"3A",X"E1",X"F0",
		X"3C",X"DD",X"BE",X"02",X"0E",X"04",X"20",X"1B",X"3A",X"E2",X"F0",X"DD",X"96",X"03",X"28",X"18",
		X"CB",X"7F",X"28",X"02",X"ED",X"44",X"FE",X"04",X"38",X"02",X"3E",X"04",X"4F",X"3A",X"E2",X"F0",
		X"DD",X"BE",X"03",X"79",X"30",X"02",X"ED",X"44",X"DD",X"77",X"06",X"3A",X"E3",X"F0",X"3C",X"DD",
		X"BE",X"04",X"3E",X"00",X"20",X"16",X"3A",X"E0",X"F0",X"DD",X"77",X"07",X"3A",X"E4",X"F0",X"DD",
		X"96",X"05",X"3E",X"00",X"28",X"06",X"3E",X"FE",X"30",X"02",X"ED",X"44",X"DD",X"77",X"09",X"18",
		X"0B",X"DD",X"7E",X"07",X"B7",X"20",X"08",X"DD",X"77",X"09",X"18",X"09",X"DD",X"7E",X"07",X"DD",
		X"86",X"09",X"DD",X"77",X"07",X"21",X"82",X"F0",X"96",X"DD",X"77",X"08",X"05",X"78",X"CB",X"27",
		X"80",X"21",X"DA",X"4C",X"85",X"30",X"01",X"24",X"6F",X"E9",X"C3",X"01",X"4D",X"C3",X"49",X"4D",
		X"C3",X"A2",X"4D",X"C3",X"12",X"4E",X"C3",X"6D",X"4E",X"C3",X"52",X"4F",X"C3",X"B0",X"4F",X"C3",
		X"F2",X"4F",X"C3",X"1C",X"50",X"C3",X"5E",X"50",X"C3",X"01",X"51",X"C3",X"60",X"51",X"C3",X"D7",
		X"51",X"0E",X"30",X"CD",X"4E",X"3D",X"FD",X"21",X"58",X"F8",X"3A",X"00",X"F0",X"47",X"FD",X"77",
		X"00",X"FD",X"36",X"02",X"40",X"3A",X"01",X"F0",X"4F",X"D6",X"08",X"FD",X"77",X"03",X"FD",X"70",
		X"04",X"FD",X"36",X"06",X"18",X"79",X"C6",X"05",X"FD",X"77",X"07",X"DD",X"34",X"00",X"DD",X"36",
		X"01",X"03",X"3A",X"82",X"F0",X"DD",X"77",X"07",X"DD",X"36",X"09",X"02",X"DD",X"36",X"06",X"00",
		X"DD",X"36",X"0A",X"02",X"DD",X"36",X"0B",X"04",X"C9",X"FD",X"21",X"58",X"F8",X"FD",X"7E",X"03",
		X"DD",X"96",X"08",X"47",X"FD",X"7E",X"07",X"DD",X"96",X"08",X"4F",X"FD",X"7E",X"05",X"EE",X"20",
		X"57",X"DD",X"35",X"01",X"20",X"32",X"DD",X"36",X"01",X"03",X"DD",X"34",X"00",X"FD",X"7E",X"00",
		X"FD",X"36",X"00",X"00",X"FD",X"36",X"04",X"00",X"FD",X"21",X"C4",X"F9",X"FD",X"77",X"00",X"FD",
		X"36",X"02",X"41",X"FD",X"77",X"04",X"DD",X"77",X"03",X"DD",X"36",X"02",X"01",X"DD",X"70",X"05",
		X"DD",X"36",X"04",X"01",X"DD",X"36",X"09",X"01",X"FD",X"70",X"03",X"FD",X"71",X"07",X"FD",X"72",
		X"05",X"C9",X"FD",X"21",X"C4",X"F9",X"CD",X"56",X"52",X"38",X"33",X"DD",X"46",X"03",X"FD",X"70",
		X"00",X"DD",X"4E",X"05",X"FD",X"71",X"03",X"DD",X"35",X"01",X"28",X"12",X"FD",X"70",X"04",X"79",
		X"C6",X"0D",X"FD",X"77",X"07",X"FD",X"7E",X"05",X"EE",X"20",X"FD",X"77",X"05",X"C9",X"78",X"DD",
		X"86",X"0A",X"FD",X"77",X"04",X"79",X"DD",X"86",X"0B",X"FD",X"77",X"07",X"18",X"0C",X"FD",X"36",
		X"00",X"00",X"FD",X"36",X"04",X"00",X"DD",X"35",X"01",X"C0",X"FD",X"34",X"02",X"FD",X"36",X"06",
		X"6C",X"DD",X"34",X"0A",X"DD",X"34",X"0B",X"3A",X"E8",X"F0",X"B7",X"20",X"04",X"DD",X"36",X"09",
		X"FF",X"DD",X"34",X"00",X"DD",X"36",X"01",X"04",X"3A",X"5D",X"F3",X"B7",X"C8",X"DD",X"36",X"01",
		X"06",X"C9",X"FD",X"21",X"C4",X"F9",X"CD",X"56",X"52",X"38",X"1C",X"DD",X"46",X"03",X"FD",X"70",
		X"00",X"DD",X"4E",X"05",X"FD",X"71",X"03",X"78",X"DD",X"86",X"0A",X"FD",X"77",X"04",X"79",X"DD",
		X"86",X"0B",X"FD",X"77",X"07",X"18",X"08",X"FD",X"36",X"00",X"00",X"FD",X"36",X"04",X"00",X"DD",
		X"34",X"0A",X"DD",X"34",X"0B",X"DD",X"35",X"01",X"C0",X"FD",X"34",X"02",X"FD",X"7E",X"02",X"FE",
		X"45",X"28",X"0E",X"DD",X"36",X"01",X"04",X"3A",X"5D",X"F3",X"B7",X"C8",X"DD",X"36",X"01",X"06",
		X"C9",X"FD",X"36",X"01",X"00",X"DD",X"36",X"01",X"0C",X"DD",X"34",X"00",X"C9",X"FD",X"21",X"C4",
		X"F9",X"CD",X"56",X"52",X"38",X"1C",X"DD",X"46",X"03",X"FD",X"70",X"00",X"DD",X"4E",X"05",X"FD",
		X"71",X"03",X"78",X"DD",X"86",X"0A",X"FD",X"77",X"04",X"79",X"DD",X"86",X"0B",X"FD",X"77",X"07",
		X"18",X"08",X"FD",X"36",X"00",X"00",X"FD",X"36",X"04",X"00",X"DD",X"35",X"01",X"28",X"0F",X"DD",
		X"34",X"0A",X"DD",X"34",X"0B",X"FD",X"7E",X"01",X"EE",X"20",X"FD",X"77",X"01",X"C9",X"FD",X"36",
		X"02",X"46",X"0E",X"19",X"CD",X"4E",X"3D",X"FD",X"36",X"04",X"00",X"DD",X"36",X"09",X"00",X"DD",
		X"7E",X"06",X"CB",X"2F",X"DD",X"77",X"06",X"3A",X"5D",X"F3",X"B7",X"C2",X"49",X"4F",X"3A",X"E8",
		X"F0",X"B7",X"CA",X"49",X"4F",X"3A",X"E1",X"F0",X"3C",X"DD",X"BE",X"02",X"C2",X"49",X"4F",X"47",
		X"3A",X"E3",X"F0",X"3C",X"DD",X"BE",X"04",X"20",X"60",X"4F",X"3A",X"E2",X"F0",X"47",X"C6",X"08",
		X"DD",X"96",X"03",X"30",X"02",X"ED",X"44",X"FE",X"0C",X"30",X"4E",X"3A",X"E4",X"F0",X"D6",X"08",
		X"DD",X"96",X"05",X"30",X"02",X"ED",X"44",X"FE",X"0C",X"30",X"3E",X"AF",X"32",X"FD",X"F0",X"32",
		X"EE",X"F0",X"21",X"60",X"B9",X"CD",X"EE",X"3D",X"21",X"E8",X"F0",X"36",X"04",X"FD",X"21",X"D8",
		X"F9",X"FD",X"36",X"00",X"00",X"21",X"DB",X"F0",X"7E",X"FE",X"09",X"20",X"0A",X"3C",X"CB",X"40",
		X"28",X"02",X"D6",X"02",X"77",X"FE",X"09",X"3E",X"FF",X"38",X"02",X"ED",X"44",X"32",X"DC",X"F0",
		X"DD",X"36",X"01",X"04",X"DD",X"36",X"00",X"06",X"C9",X"DD",X"36",X"01",X"04",X"DD",X"36",X"00",
		X"0C",X"C9",X"CD",X"56",X"52",X"FD",X"21",X"C4",X"F9",X"38",X"0E",X"DD",X"7E",X"03",X"FD",X"77",
		X"00",X"DD",X"7E",X"05",X"FD",X"77",X"03",X"18",X"04",X"FD",X"36",X"00",X"00",X"DD",X"35",X"01",
		X"C0",X"21",X"DB",X"F0",X"7E",X"FE",X"09",X"28",X"12",X"3A",X"DC",X"F0",X"86",X"CB",X"7F",X"20",
		X"07",X"FE",X"0C",X"38",X"05",X"AF",X"18",X"02",X"3E",X"0B",X"77",X"FD",X"7E",X"02",X"3C",X"FE",
		X"4B",X"28",X"10",X"FD",X"77",X"02",X"DD",X"36",X"01",X"04",X"7E",X"FE",X"09",X"C0",X"DD",X"36",
		X"00",X"07",X"C9",X"FD",X"36",X"00",X"00",X"DD",X"36",X"00",X"08",X"DD",X"36",X"01",X"04",X"C9",
		X"CD",X"56",X"52",X"FD",X"21",X"C4",X"F9",X"38",X"0E",X"DD",X"7E",X"03",X"FD",X"77",X"00",X"DD",
		X"7E",X"05",X"FD",X"77",X"03",X"18",X"04",X"FD",X"36",X"00",X"00",X"DD",X"35",X"01",X"C0",X"FD",
		X"7E",X"02",X"3C",X"FE",X"4B",X"28",X"09",X"FD",X"77",X"02",X"DD",X"36",X"00",X"09",X"18",X"08",
		X"FD",X"36",X"00",X"00",X"DD",X"36",X"00",X"0A",X"DD",X"36",X"01",X"04",X"21",X"DB",X"F0",X"36",
		X"0C",X"C9",X"DD",X"35",X"01",X"C0",X"DD",X"36",X"01",X"04",X"21",X"DB",X"F0",X"7E",X"FE",X"09",
		X"28",X"13",X"3A",X"DC",X"F0",X"86",X"CB",X"7F",X"20",X"07",X"FE",X"0C",X"38",X"05",X"AF",X"18",
		X"02",X"3E",X"0B",X"77",X"C9",X"36",X"0C",X"DD",X"36",X"00",X"0A",X"C9",X"CD",X"56",X"52",X"FD",
		X"21",X"C4",X"F9",X"38",X"0E",X"DD",X"7E",X"03",X"FD",X"77",X"00",X"DD",X"7E",X"05",X"FD",X"77",
		X"03",X"18",X"04",X"FD",X"36",X"00",X"00",X"DD",X"35",X"01",X"C0",X"DD",X"36",X"01",X"06",X"FD",
		X"7E",X"02",X"3C",X"FE",X"4B",X"28",X"05",X"FD",X"77",X"02",X"18",X"08",X"FD",X"36",X"00",X"00",
		X"DD",X"36",X"00",X"0B",X"3A",X"DB",X"F0",X"FE",X"09",X"20",X"0E",X"C3",X"05",X"51",X"DD",X"35",
		X"01",X"C0",X"DD",X"36",X"01",X"06",X"DD",X"34",X"00",X"AF",X"32",X"D9",X"F0",X"32",X"E8",X"F0",
		X"21",X"DB",X"F0",X"36",X"09",X"0E",X"15",X"CD",X"4E",X"3D",X"11",X"04",X"00",X"FD",X"21",X"CC",
		X"F9",X"FD",X"36",X"00",X"00",X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",X"19",X"FD",X"36",X"00",
		X"00",X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",X"19",X"CD",X"43",X"51",X"CD",X"13",X"5C",X"11",
		X"04",X"00",X"FD",X"21",X"DC",X"F9",X"FD",X"36",X"02",X"52",X"FD",X"36",X"01",X"00",X"3A",X"E2",
		X"F0",X"47",X"D6",X"10",X"6F",X"3A",X"E4",X"F0",X"4F",X"D6",X"10",X"CB",X"4C",X"28",X"06",X"FD",
		X"70",X"00",X"FD",X"77",X"03",X"FD",X"19",X"CB",X"54",X"28",X"0E",X"FD",X"70",X"00",X"FD",X"36",
		X"02",X"53",X"FD",X"36",X"01",X"00",X"FD",X"71",X"03",X"FD",X"19",X"CB",X"44",X"28",X"0E",X"FD",
		X"75",X"00",X"FD",X"36",X"02",X"54",X"FD",X"36",X"01",X"00",X"FD",X"77",X"03",X"FD",X"19",X"CB",
		X"5C",X"C8",X"FD",X"75",X"00",X"FD",X"36",X"02",X"55",X"FD",X"36",X"01",X"00",X"FD",X"71",X"03",
		X"C9",X"DD",X"35",X"01",X"C0",X"11",X"04",X"00",X"FD",X"21",X"DC",X"F9",X"FD",X"7E",X"02",X"C6",
		X"04",X"FE",X"5E",X"28",X"26",X"FD",X"77",X"02",X"FD",X"19",X"FD",X"7E",X"02",X"C6",X"04",X"FD",
		X"77",X"02",X"FD",X"19",X"FD",X"7E",X"02",X"C6",X"04",X"FD",X"77",X"02",X"FD",X"19",X"FD",X"7E",
		X"02",X"C6",X"04",X"FD",X"77",X"02",X"DD",X"36",X"01",X"06",X"C9",X"DD",X"36",X"00",X"0D",X"DD",
		X"36",X"01",X"10",X"FD",X"36",X"00",X"00",X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",X"19",X"FD",
		X"36",X"00",X"00",X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",X"19",X"FD",X"36",X"00",X"00",X"C9",
		X"3A",X"5D",X"F3",X"B7",X"CC",X"56",X"52",X"FD",X"21",X"C4",X"F9",X"38",X"0E",X"DD",X"7E",X"03",
		X"FD",X"77",X"00",X"DD",X"7E",X"05",X"FD",X"77",X"03",X"18",X"04",X"FD",X"36",X"00",X"00",X"DD",
		X"35",X"01",X"C0",X"FD",X"7E",X"02",X"3C",X"FE",X"4B",X"28",X"08",X"FD",X"77",X"02",X"DD",X"36",
		X"01",X"04",X"C9",X"FD",X"36",X"00",X"00",X"DD",X"36",X"00",X"0D",X"DD",X"36",X"01",X"10",X"3A",
		X"5D",X"F3",X"B7",X"C8",X"DD",X"36",X"00",X"00",X"2A",X"9B",X"F0",X"3A",X"68",X"F3",X"FE",X"1A",
		X"30",X"1B",X"C6",X"41",X"77",X"7D",X"FE",X"8C",X"20",X"05",X"3E",X"02",X"32",X"6B",X"F3",X"2B",
		X"2B",X"22",X"9B",X"F0",X"3A",X"E2",X"F0",X"C6",X"10",X"32",X"E2",X"F0",X"C9",X"20",X"03",X"36",
		X"00",X"C9",X"AF",X"32",X"E8",X"F0",X"C9",X"DD",X"35",X"01",X"C0",X"0E",X"1A",X"CD",X"4E",X"3D",
		X"3A",X"E8",X"F0",X"B7",X"28",X"05",X"0E",X"2B",X"CD",X"4E",X"3D",X"DD",X"36",X"00",X"00",X"C9",
		X"21",X"FE",X"F0",X"7E",X"B7",X"20",X"0E",X"3A",X"12",X"F0",X"47",X"E6",X"80",X"C8",X"78",X"EE",
		X"80",X"32",X"12",X"F0",X"C9",X"3A",X"03",X"F0",X"E6",X"13",X"C0",X"DB",X"01",X"2F",X"E6",X"02",
		X"C8",X"35",X"DD",X"34",X"00",X"3A",X"5D",X"F3",X"B7",X"C8",X"AF",X"32",X"6D",X"F3",X"3A",X"68",
		X"F3",X"FE",X"0E",X"3E",X"02",X"30",X"01",X"AF",X"32",X"E0",X"F0",X"3A",X"68",X"F3",X"D6",X"1A",
		X"38",X"1A",X"C0",X"32",X"6B",X"F3",X"2A",X"9B",X"F0",X"7D",X"FE",X"90",X"28",X"13",X"23",X"23",
		X"22",X"9B",X"F0",X"3A",X"E2",X"F0",X"D6",X"10",X"32",X"E2",X"F0",X"C9",X"3A",X"6B",X"F3",X"B7",
		X"C8",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"7E",X"06",X"B7",X"28",X"19",X"CB",X"7F",X"20",X"0A",
		X"DD",X"86",X"03",X"30",X"0D",X"DD",X"34",X"02",X"18",X"08",X"DD",X"86",X"03",X"38",X"03",X"DD",
		X"35",X"02",X"DD",X"77",X"03",X"DD",X"7E",X"08",X"ED",X"44",X"28",X"19",X"CB",X"7F",X"20",X"0A",
		X"DD",X"86",X"05",X"30",X"0D",X"DD",X"34",X"04",X"18",X"08",X"DD",X"86",X"05",X"38",X"03",X"DD",
		X"35",X"04",X"DD",X"77",X"05",X"DD",X"7E",X"02",X"DD",X"A6",X"04",X"FE",X"01",X"C8",X"37",X"C9",
		X"3A",X"D2",X"F0",X"B7",X"20",X"0E",X"3A",X"12",X"F0",X"47",X"E6",X"08",X"C8",X"78",X"EE",X"08",
		X"32",X"12",X"F0",X"C9",X"3A",X"03",X"F0",X"47",X"E6",X"10",X"20",X"12",X"78",X"E6",X"03",X"28",
		X"06",X"AF",X"32",X"D2",X"F0",X"18",X"07",X"DB",X"01",X"2F",X"E6",X"01",X"20",X"08",X"3A",X"D3",
		X"F0",X"B7",X"C8",X"C3",X"F5",X"53",X"3A",X"D3",X"F0",X"B7",X"20",X"09",X"0E",X"24",X"CD",X"4E",
		X"3D",X"3C",X"32",X"D3",X"F0",X"3A",X"15",X"F0",X"B7",X"C2",X"8E",X"53",X"FD",X"21",X"54",X"F8",
		X"3A",X"00",X"F0",X"FD",X"77",X"00",X"47",X"3A",X"01",X"F0",X"4F",X"C6",X"14",X"FD",X"77",X"03",
		X"FD",X"7E",X"01",X"EE",X"20",X"FD",X"77",X"01",X"FD",X"36",X"02",X"15",X"3A",X"FF",X"F0",X"B7",
		X"28",X"04",X"FE",X"03",X"38",X"26",X"FD",X"21",X"58",X"F8",X"78",X"D6",X"04",X"FD",X"77",X"00",
		X"79",X"C6",X"1C",X"FD",X"77",X"03",X"FD",X"36",X"02",X"2E",X"11",X"04",X"00",X"FD",X"19",X"FD",
		X"77",X"03",X"78",X"C6",X"04",X"FD",X"77",X"00",X"FD",X"36",X"02",X"2E",X"2A",X"81",X"F0",X"ED",
		X"5B",X"D0",X"F0",X"19",X"7C",X"D6",X"0C",X"30",X"04",X"22",X"D0",X"F0",X"C9",X"67",X"22",X"D0",
		X"F0",X"81",X"57",X"CD",X"B3",X"3D",X"CD",X"E4",X"3D",X"78",X"D6",X"04",X"FD",X"77",X"00",X"7A",
		X"C6",X"1C",X"FD",X"77",X"03",X"FD",X"36",X"02",X"2E",X"36",X"03",X"CD",X"B3",X"3D",X"CD",X"E4",
		X"3D",X"78",X"C6",X"04",X"FD",X"77",X"00",X"7A",X"C6",X"1C",X"FD",X"77",X"03",X"FD",X"36",X"02",
		X"2E",X"36",X"03",X"21",X"D2",X"F0",X"35",X"28",X"6C",X"2A",X"D0",X"F0",X"18",X"B6",X"21",X"00",
		X"F0",X"46",X"23",X"4E",X"2A",X"81",X"F0",X"ED",X"5B",X"D0",X"F0",X"19",X"7C",X"D6",X"08",X"30",
		X"04",X"22",X"D0",X"F0",X"C9",X"67",X"22",X"D0",X"F0",X"81",X"57",X"3A",X"D2",X"F0",X"E6",X"03",
		X"5F",X"CD",X"B3",X"3D",X"CD",X"E4",X"3D",X"78",X"D6",X"03",X"93",X"FD",X"77",X"00",X"7A",X"C6",
		X"1C",X"FD",X"77",X"03",X"3E",X"9C",X"83",X"FD",X"77",X"02",X"36",X"28",X"CD",X"B3",X"3D",X"CD",
		X"E4",X"3D",X"78",X"C6",X"09",X"93",X"FD",X"77",X"00",X"7A",X"C6",X"1C",X"FD",X"77",X"03",X"7B",
		X"3C",X"E6",X"03",X"C6",X"9C",X"FD",X"77",X"02",X"36",X"28",X"21",X"D2",X"F0",X"35",X"28",X"05",
		X"2A",X"D0",X"F0",X"18",X"A7",X"0E",X"21",X"CD",X"4E",X"3D",X"AF",X"32",X"D3",X"F0",X"32",X"D0",
		X"F0",X"32",X"D1",X"F0",X"3A",X"15",X"F0",X"B7",X"C0",X"32",X"54",X"F8",X"3A",X"FF",X"F0",X"B7",
		X"28",X"04",X"FE",X"03",X"D8",X"AF",X"32",X"58",X"F8",X"32",X"5C",X"F8",X"C9",X"3A",X"D8",X"F0",
		X"B7",X"CA",X"A1",X"54",X"47",X"DD",X"21",X"00",X"F9",X"21",X"0B",X"F1",X"0E",X"F0",X"3A",X"01",
		X"F0",X"FE",X"90",X"30",X"03",X"C6",X"60",X"4F",X"DD",X"7E",X"00",X"B7",X"28",X"59",X"DD",X"7E",
		X"03",X"C6",X"0C",X"B9",X"38",X"22",X"DD",X"7E",X"02",X"FE",X"19",X"28",X"0E",X"DD",X"36",X"02",
		X"19",X"DD",X"7E",X"03",X"C6",X"04",X"DD",X"77",X"03",X"18",X"3B",X"DD",X"36",X"00",X"00",X"3A",
		X"D8",X"F0",X"3D",X"32",X"D8",X"F0",X"18",X"2E",X"DD",X"77",X"03",X"7E",X"B7",X"28",X"27",X"57",
		X"DD",X"86",X"00",X"FE",X"08",X"38",X"19",X"FE",X"F8",X"30",X"15",X"5F",X"CD",X"98",X"3F",X"E5",
		X"CD",X"DA",X"3F",X"FD",X"73",X"00",X"72",X"E1",X"DD",X"7E",X"03",X"D6",X"02",X"FD",X"77",X"03",
		X"36",X"00",X"DD",X"36",X"02",X"2F",X"05",X"11",X"04",X"00",X"DD",X"19",X"23",X"78",X"B7",X"20",
		X"97",X"3A",X"D5",X"F0",X"B7",X"CA",X"5C",X"55",X"3A",X"03",X"F0",X"E6",X"13",X"28",X"07",X"AF",
		X"32",X"D5",X"F0",X"C3",X"52",X"55",X"3A",X"D7",X"F0",X"B7",X"28",X"05",X"3D",X"32",X"D7",X"F0",
		X"C9",X"3A",X"D6",X"F0",X"B7",X"20",X"1B",X"3C",X"32",X"D6",X"F0",X"FD",X"21",X"FC",X"F8",X"FD",
		X"36",X"00",X"00",X"FD",X"36",X"02",X"18",X"0E",X"25",X"CD",X"4E",X"3D",X"21",X"24",X"F0",X"36",
		X"04",X"C9",X"4F",X"FD",X"21",X"FC",X"F8",X"3A",X"00",X"F0",X"57",X"FD",X"77",X"00",X"3A",X"01",
		X"F0",X"5F",X"C6",X"14",X"FD",X"77",X"03",X"FD",X"7E",X"01",X"EE",X"20",X"FD",X"77",X"01",X"0D",
		X"20",X"0A",X"21",X"D6",X"F0",X"34",X"21",X"D7",X"F0",X"36",X"02",X"C9",X"CD",X"98",X"3F",X"CD",
		X"DA",X"3F",X"7A",X"C6",X"06",X"FD",X"77",X"00",X"7B",X"C6",X"1C",X"FD",X"77",X"03",X"CB",X"47",
		X"28",X"08",X"FD",X"7E",X"01",X"EE",X"10",X"FD",X"77",X"01",X"36",X"06",X"CD",X"98",X"3F",X"CD",
		X"DA",X"3F",X"7A",X"D6",X"06",X"FD",X"77",X"00",X"7B",X"C6",X"1A",X"FD",X"77",X"03",X"CB",X"7F",
		X"20",X"08",X"FD",X"7E",X"01",X"EE",X"10",X"FD",X"77",X"01",X"36",X"FA",X"21",X"D5",X"F0",X"35",
		X"C0",X"AF",X"32",X"FC",X"F8",X"32",X"D0",X"F0",X"32",X"D6",X"F0",X"C9",X"3A",X"03",X"F0",X"E6",
		X"10",X"C0",X"21",X"D4",X"F0",X"7E",X"B7",X"28",X"0D",X"DB",X"01",X"2F",X"E6",X"08",X"C8",X"35",
		X"21",X"D5",X"F0",X"36",X"40",X"C9",X"3A",X"12",X"F0",X"E6",X"02",X"C8",X"3A",X"12",X"F0",X"EE",
		X"02",X"32",X"12",X"F0",X"C9",X"3A",X"15",X"F0",X"B7",X"20",X"33",X"06",X"02",X"11",X"04",X"00",
		X"DD",X"21",X"60",X"F8",X"21",X"53",X"F0",X"DD",X"7E",X"00",X"B7",X"28",X"1D",X"86",X"FE",X"10",
		X"38",X"0E",X"DD",X"77",X"00",X"3A",X"52",X"F0",X"DD",X"86",X"03",X"DD",X"77",X"03",X"18",X"0E",
		X"DD",X"36",X"00",X"00",X"DD",X"36",X"03",X"00",X"18",X"04",X"DD",X"19",X"10",X"D9",X"3A",X"43",
		X"F0",X"FE",X"01",X"38",X"1E",X"CA",X"4F",X"58",X"3D",X"32",X"43",X"F0",X"FE",X"01",X"20",X"13",
		X"3A",X"49",X"F0",X"B7",X"28",X"07",X"3E",X"02",X"32",X"43",X"F0",X"18",X"06",X"32",X"44",X"F0",
		X"32",X"2F",X"F0",X"3A",X"46",X"F0",X"B7",X"C8",X"DD",X"2A",X"48",X"F0",X"DD",X"7E",X"08",X"B7",
		X"C0",X"3A",X"03",X"F0",X"E6",X"13",X"28",X"17",X"21",X"46",X"F0",X"36",X"00",X"DD",X"36",X"0D",
		X"01",X"AF",X"32",X"4B",X"F0",X"32",X"4C",X"F0",X"32",X"55",X"F1",X"32",X"D8",X"F8",X"C9",X"DD",
		X"7E",X"01",X"47",X"E6",X"0A",X"20",X"E1",X"78",X"E6",X"04",X"20",X"E1",X"FD",X"21",X"D8",X"F8",
		X"FD",X"7E",X"00",X"B7",X"28",X"1C",X"DD",X"7E",X"07",X"FE",X"11",X"38",X"D0",X"FE",X"E0",X"30",
		X"CC",X"DD",X"7E",X"07",X"C6",X"10",X"FD",X"77",X"03",X"3A",X"55",X"F1",X"DD",X"86",X"05",X"FD",
		X"77",X"00",X"3A",X"42",X"F0",X"B7",X"20",X"0B",X"3A",X"4C",X"F0",X"B7",X"28",X"05",X"3D",X"32",
		X"4C",X"F0",X"C9",X"3A",X"4A",X"F0",X"B7",X"20",X"3B",X"3A",X"00",X"F0",X"DD",X"96",X"05",X"30",
		X"02",X"ED",X"44",X"D6",X"08",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"B7",X"47",X"3A",
		X"01",X"F0",X"28",X"05",X"DD",X"96",X"10",X"10",X"FB",X"D6",X"08",X"DD",X"BE",X"07",X"D8",X"D6",
		X"08",X"DD",X"BE",X"07",X"D0",X"3A",X"42",X"F0",X"B7",X"20",X"09",X"3A",X"06",X"F0",X"DD",X"BE",
		X"09",X"C2",X"F8",X"55",X"3A",X"4B",X"F0",X"47",X"CB",X"27",X"80",X"21",X"A4",X"56",X"85",X"30",
		X"01",X"24",X"6F",X"E9",X"C3",X"B3",X"56",X"C3",X"EE",X"56",X"C3",X"36",X"57",X"C3",X"C2",X"57",
		X"C3",X"0C",X"58",X"21",X"00",X"F0",X"DD",X"7E",X"05",X"BE",X"38",X"0D",X"D6",X"0C",X"FD",X"77",
		X"00",X"FD",X"36",X"01",X"20",X"3E",X"F4",X"18",X"0B",X"C6",X"0C",X"FD",X"77",X"00",X"FD",X"36",
		X"01",X"00",X"3E",X"0C",X"32",X"55",X"F1",X"FD",X"36",X"02",X"10",X"DD",X"7E",X"07",X"C6",X"10",
		X"FD",X"77",X"03",X"3A",X"4D",X"F0",X"32",X"4C",X"F0",X"21",X"4B",X"F0",X"34",X"C9",X"21",X"00",
		X"F0",X"DD",X"7E",X"05",X"BE",X"3E",X"0C",X"38",X"02",X"ED",X"44",X"21",X"55",X"F1",X"BE",X"20",
		X"1A",X"0E",X"11",X"CD",X"4E",X"3D",X"21",X"4E",X"F0",X"36",X"02",X"3A",X"4D",X"F0",X"32",X"4C",
		X"F0",X"21",X"4B",X"F0",X"34",X"21",X"4A",X"F0",X"36",X"00",X"C9",X"21",X"4B",X"F0",X"36",X"00",
		X"21",X"4C",X"F0",X"36",X"10",X"FD",X"36",X"00",X"00",X"FD",X"36",X"02",X"00",X"FD",X"36",X"03",
		X"00",X"FD",X"36",X"01",X"00",X"C9",X"21",X"00",X"F0",X"DD",X"7E",X"05",X"BE",X"57",X"5E",X"3E",
		X"0C",X"38",X"04",X"ED",X"44",X"5A",X"56",X"21",X"55",X"F1",X"BE",X"20",X"CE",X"3A",X"42",X"F0",
		X"B7",X"20",X"47",X"DD",X"7E",X"07",X"C6",X"14",X"47",X"0E",X"00",X"DD",X"21",X"8B",X"F2",X"79",
		X"FE",X"06",X"28",X"3C",X"DD",X"7E",X"01",X"E6",X"80",X"28",X"25",X"DD",X"7E",X"02",X"E6",X"0F",
		X"28",X"1E",X"DD",X"7E",X"08",X"B7",X"20",X"18",X"78",X"DD",X"BE",X"07",X"38",X"12",X"DD",X"96",
		X"0E",X"D6",X"04",X"DD",X"BE",X"07",X"30",X"08",X"DD",X"7E",X"05",X"BA",X"38",X"02",X"BB",X"D8",
		X"D5",X"11",X"23",X"00",X"DD",X"19",X"D1",X"0C",X"18",X"C5",X"3A",X"82",X"F0",X"FE",X"0E",X"D0",
		X"FD",X"7E",X"02",X"3C",X"FD",X"77",X"02",X"0E",X"1B",X"CD",X"4E",X"3D",X"FD",X"7E",X"00",X"32",
		X"4F",X"F0",X"FD",X"7E",X"03",X"32",X"50",X"F0",X"21",X"4B",X"F0",X"34",X"21",X"4A",X"F0",X"36",
		X"01",X"C9",X"3A",X"55",X"F1",X"B7",X"3E",X"10",X"06",X"00",X"F2",X"D1",X"57",X"ED",X"44",X"06",
		X"20",X"4F",X"DD",X"7E",X"10",X"32",X"52",X"F0",X"3A",X"4E",X"F0",X"3D",X"DD",X"21",X"60",X"F8",
		X"21",X"53",X"F0",X"28",X"04",X"DD",X"21",X"64",X"F8",X"DD",X"70",X"01",X"DD",X"36",X"02",X"12",
		X"71",X"3A",X"50",X"F0",X"21",X"52",X"F0",X"86",X"DD",X"77",X"03",X"3A",X"4F",X"F0",X"81",X"DD",
		X"77",X"00",X"21",X"4C",X"F0",X"36",X"08",X"21",X"4B",X"F0",X"34",X"C9",X"0E",X"1C",X"CD",X"4E",
		X"3D",X"FD",X"7E",X"02",X"3D",X"FD",X"77",X"02",X"21",X"4A",X"F0",X"36",X"00",X"3A",X"4E",X"F0",
		X"3D",X"32",X"4E",X"F0",X"20",X"1B",X"21",X"4B",X"F0",X"36",X"00",X"21",X"4C",X"F0",X"36",X"20",
		X"FD",X"36",X"00",X"00",X"FD",X"36",X"02",X"00",X"FD",X"36",X"03",X"00",X"FD",X"36",X"01",X"00",
		X"C9",X"21",X"4B",X"F0",X"36",X"02",X"3A",X"4D",X"F0",X"CB",X"27",X"32",X"4C",X"F0",X"C9",X"3A",
		X"15",X"F0",X"B7",X"20",X"06",X"3A",X"33",X"F0",X"B7",X"20",X"16",X"21",X"E7",X"F0",X"36",X"02",
		X"3A",X"E5",X"F0",X"B7",X"C2",X"18",X"5A",X"3C",X"32",X"E5",X"F0",X"32",X"E6",X"F0",X"C3",X"18",
		X"5A",X"3A",X"44",X"F0",X"47",X"CB",X"27",X"80",X"21",X"81",X"58",X"85",X"30",X"01",X"24",X"6F",
		X"E9",X"C3",X"8A",X"58",X"C3",X"4E",X"59",X"C3",X"DB",X"59",X"3A",X"06",X"F0",X"FE",X"02",X"30",
		X"0D",X"3A",X"09",X"F0",X"B7",X"20",X"07",X"3A",X"82",X"F0",X"B7",X"C2",X"18",X"5A",X"DD",X"21",
		X"8B",X"F2",X"06",X"06",X"11",X"23",X"00",X"DD",X"7E",X"01",X"B7",X"28",X"1B",X"DD",X"19",X"10",
		X"F6",X"DD",X"21",X"8B",X"F2",X"06",X"06",X"DD",X"7E",X"05",X"B7",X"28",X"08",X"DD",X"19",X"10",
		X"F6",X"DD",X"21",X"8B",X"F2",X"CD",X"32",X"3F",X"21",X"32",X"F0",X"34",X"DD",X"22",X"48",X"F0",
		X"06",X"00",X"0E",X"F7",X"FD",X"21",X"5B",X"F2",X"CD",X"B5",X"41",X"21",X"00",X"F0",X"FD",X"7E",
		X"02",X"B7",X"28",X"03",X"BE",X"38",X"03",X"FD",X"7E",X"00",X"D6",X"10",X"30",X"08",X"FD",X"7E",
		X"02",X"D6",X"10",X"DA",X"18",X"5A",X"DD",X"77",X"05",X"DD",X"36",X"07",X"F7",X"DD",X"36",X"08",
		X"00",X"DD",X"36",X"01",X"83",X"3A",X"82",X"F0",X"DD",X"77",X"03",X"DD",X"36",X"0B",X"0C",X"DD",
		X"36",X"04",X"00",X"DD",X"36",X"02",X"10",X"DD",X"36",X"06",X"25",X"DD",X"36",X"1D",X"26",X"DD",
		X"36",X"1E",X"00",X"3A",X"E1",X"BA",X"DD",X"77",X"0E",X"3A",X"EA",X"BA",X"DD",X"77",X"0F",X"3A",
		X"06",X"F0",X"DD",X"77",X"09",X"DD",X"36",X"1F",X"00",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"10",
		X"00",X"3E",X"01",X"32",X"46",X"F0",X"32",X"44",X"F0",X"AF",X"32",X"42",X"F0",X"C9",X"DD",X"2A",
		X"48",X"F0",X"3A",X"82",X"F0",X"DD",X"77",X"03",X"3A",X"06",X"F0",X"FE",X"02",X"38",X"72",X"DD",
		X"77",X"09",X"3A",X"01",X"F0",X"D6",X"0A",X"DD",X"BE",X"07",X"3E",X"00",X"28",X"06",X"38",X"03",
		X"3D",X"18",X"01",X"3C",X"DD",X"77",X"10",X"ED",X"44",X"DD",X"86",X"07",X"DD",X"77",X"07",X"4F",
		X"06",X"00",X"FD",X"21",X"5B",X"F2",X"CD",X"B5",X"41",X"21",X"00",X"F0",X"FD",X"7E",X"02",X"B7",
		X"28",X"03",X"BE",X"38",X"03",X"FD",X"7E",X"00",X"D6",X"10",X"30",X"05",X"FD",X"7E",X"02",X"D6",
		X"10",X"47",X"DD",X"96",X"05",X"30",X"02",X"ED",X"44",X"FE",X"10",X"38",X"0A",X"DD",X"36",X"03",
		X"00",X"21",X"43",X"F0",X"36",X"20",X"C9",X"DD",X"70",X"05",X"DD",X"36",X"01",X"80",X"CD",X"E3",
		X"55",X"DD",X"2A",X"48",X"F0",X"DD",X"36",X"01",X"83",X"3A",X"03",X"F0",X"E6",X"02",X"20",X"06",
		X"C9",X"21",X"42",X"F0",X"36",X"01",X"21",X"44",X"F0",X"34",X"C9",X"DD",X"2A",X"48",X"F0",X"DD",
		X"36",X"01",X"80",X"DD",X"7E",X"05",X"C6",X"04",X"DD",X"77",X"05",X"DD",X"36",X"0B",X"02",X"DD",
		X"36",X"03",X"01",X"DD",X"36",X"0D",X"40",X"3A",X"09",X"F0",X"B7",X"28",X"09",X"3A",X"82",X"F0",
		X"3C",X"DD",X"77",X"03",X"18",X"06",X"3A",X"82",X"F0",X"B7",X"20",X"04",X"DD",X"36",X"0B",X"0C",
		X"DD",X"36",X"04",X"02",X"DD",X"36",X"0C",X"04",X"21",X"43",X"F0",X"36",X"00",X"C9",X"3A",X"D9",
		X"F0",X"FE",X"01",X"D8",X"20",X"04",X"3C",X"32",X"D9",X"F0",X"21",X"E2",X"F0",X"46",X"21",X"E4",
		X"F0",X"4E",X"21",X"71",X"BB",X"3A",X"DB",X"F0",X"CB",X"27",X"57",X"CB",X"27",X"CB",X"27",X"82",
		X"85",X"30",X"01",X"24",X"6F",X"E5",X"FD",X"E1",X"CD",X"13",X"5C",X"11",X"04",X"00",X"DD",X"21",
		X"CC",X"F9",X"7C",X"E6",X"80",X"28",X"0F",X"FD",X"7E",X"09",X"DD",X"77",X"02",X"79",X"C6",X"04",
		X"DD",X"77",X"03",X"78",X"C6",X"14",X"DD",X"77",X"00",X"DD",X"21",X"D0",X"F9",X"7C",X"E6",X"10",
		X"28",X"17",X"FD",X"7E",X"01",X"DD",X"77",X"02",X"FD",X"7E",X"04",X"DD",X"77",X"01",X"FD",X"7E",
		X"02",X"81",X"DD",X"77",X"03",X"FD",X"7E",X"00",X"80",X"DD",X"77",X"00",X"DD",X"19",X"7C",X"E6",
		X"20",X"28",X"1E",X"FD",X"7E",X"01",X"FE",X"51",X"20",X"02",X"3E",X"03",X"3C",X"DD",X"77",X"02",
		X"FD",X"7E",X"04",X"DD",X"77",X"01",X"FD",X"7E",X"05",X"81",X"DD",X"77",X"03",X"FD",X"7E",X"03",
		X"80",X"DD",X"77",X"00",X"DD",X"21",X"DC",X"F9",X"3A",X"D9",X"F0",X"FE",X"02",X"3A",X"DA",X"F0",
		X"C2",X"69",X"5B",X"CB",X"4F",X"28",X"76",X"CB",X"44",X"28",X"11",X"DD",X"70",X"00",X"DD",X"36",
		X"02",X"0B",X"DD",X"36",X"01",X"20",X"79",X"D6",X"10",X"DD",X"77",X"03",X"CB",X"4C",X"28",X"16",
		X"DD",X"19",X"78",X"C6",X"10",X"DD",X"77",X"00",X"DD",X"36",X"02",X"0B",X"DD",X"36",X"01",X"00",
		X"79",X"D6",X"10",X"DD",X"77",X"03",X"CB",X"54",X"28",X"13",X"DD",X"19",X"78",X"C6",X"10",X"DD",
		X"77",X"00",X"DD",X"36",X"02",X"0B",X"DD",X"36",X"01",X"10",X"DD",X"71",X"03",X"CB",X"5C",X"28",
		X"10",X"DD",X"19",X"DD",X"70",X"00",X"DD",X"36",X"02",X"0B",X"DD",X"36",X"01",X"30",X"DD",X"71",
		X"03",X"CB",X"74",X"28",X"34",X"DD",X"19",X"FD",X"7E",X"06",X"80",X"DD",X"77",X"00",X"FD",X"7E",
		X"07",X"DD",X"77",X"02",X"FD",X"7E",X"08",X"81",X"DD",X"77",X"03",X"18",X"1C",X"DD",X"36",X"00",
		X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",X"19",X"DD",
		X"36",X"00",X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"21",X"DA",X"F0",X"7E",X"B7",X"20",X"07",
		X"36",X"0C",X"21",X"D9",X"F0",X"34",X"C9",X"35",X"C9",X"CB",X"4F",X"28",X"7C",X"CB",X"44",X"28",
		X"11",X"DD",X"70",X"00",X"DD",X"36",X"02",X"0C",X"DD",X"36",X"01",X"20",X"79",X"D6",X"10",X"DD",
		X"77",X"03",X"CB",X"4C",X"28",X"16",X"DD",X"19",X"78",X"C6",X"10",X"DD",X"77",X"00",X"DD",X"36",
		X"02",X"0C",X"DD",X"36",X"01",X"00",X"79",X"D6",X"10",X"DD",X"77",X"03",X"CB",X"54",X"28",X"13",
		X"DD",X"19",X"78",X"C6",X"10",X"DD",X"77",X"00",X"DD",X"36",X"02",X"0C",X"DD",X"36",X"01",X"10",
		X"DD",X"71",X"03",X"CB",X"5C",X"28",X"10",X"DD",X"19",X"DD",X"70",X"00",X"DD",X"36",X"02",X"0C",
		X"DD",X"36",X"01",X"30",X"DD",X"71",X"03",X"CB",X"74",X"28",X"3A",X"DD",X"19",X"FD",X"7E",X"06",
		X"80",X"DD",X"77",X"00",X"FD",X"7E",X"07",X"DD",X"77",X"02",X"FD",X"7E",X"04",X"DD",X"77",X"01",
		X"FD",X"7E",X"08",X"81",X"DD",X"77",X"03",X"18",X"1C",X"DD",X"36",X"00",X"00",X"DD",X"19",X"DD",
		X"36",X"00",X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",
		X"19",X"DD",X"36",X"00",X"00",X"21",X"DA",X"F0",X"7E",X"B7",X"20",X"05",X"36",X"0C",X"21",X"D9",
		X"F0",X"35",X"C9",X"3A",X"DB",X"F0",X"57",X"CB",X"27",X"82",X"57",X"21",X"24",X"5C",X"85",X"30",
		X"01",X"24",X"6F",X"E9",X"C3",X"48",X"5C",X"C3",X"7D",X"5C",X"C3",X"C0",X"5C",X"C3",X"C0",X"5C",
		X"C3",X"C0",X"5C",X"C3",X"7D",X"5C",X"C3",X"48",X"5C",X"C3",X"48",X"5C",X"C3",X"FA",X"5C",X"C3",
		X"FA",X"5C",X"C3",X"FA",X"5C",X"C3",X"48",X"5C",X"3A",X"E3",X"F0",X"FE",X"01",X"79",X"28",X"21",
		X"38",X"0C",X"1E",X"00",X"FE",X"FC",X"DA",X"40",X"5D",X"1E",X"8C",X"C3",X"40",X"5D",X"1E",X"FC",
		X"FE",X"09",X"DA",X"40",X"5D",X"1E",X"FF",X"FE",X"F9",X"DA",X"40",X"5D",X"1E",X"73",X"C3",X"40",
		X"5D",X"1E",X"03",X"FE",X"09",X"DA",X"40",X"5D",X"1E",X"00",X"C3",X"40",X"5D",X"3A",X"E3",X"F0",
		X"FE",X"01",X"79",X"28",X"28",X"38",X"0C",X"1E",X"00",X"FE",X"FA",X"DA",X"40",X"5D",X"1E",X"0C",
		X"C3",X"40",X"5D",X"1E",X"9C",X"FE",X"05",X"DA",X"40",X"5D",X"1E",X"BC",X"FE",X"09",X"DA",X"40",
		X"5D",X"1E",X"FF",X"FE",X"F7",X"DA",X"40",X"5D",X"1E",X"73",X"C3",X"40",X"5D",X"1E",X"73",X"FE",
		X"04",X"DA",X"40",X"5D",X"1E",X"43",X"FE",X"09",X"DA",X"40",X"5D",X"1E",X"00",X"C3",X"40",X"5D",
		X"3A",X"E3",X"F0",X"FE",X"01",X"79",X"28",X"22",X"38",X"0A",X"1E",X"00",X"FE",X"F9",X"38",X"70",
		X"1E",X"8C",X"18",X"6C",X"1E",X"9C",X"FE",X"09",X"38",X"66",X"1E",X"9F",X"FE",X"11",X"38",X"60",
		X"1E",X"FF",X"FE",X"F9",X"38",X"5A",X"1E",X"73",X"18",X"56",X"1E",X"63",X"FE",X"09",X"38",X"50",
		X"1E",X"60",X"FE",X"10",X"38",X"4A",X"1E",X"00",X"18",X"46",X"3A",X"E3",X"F0",X"FE",X"01",X"79",
		X"28",X"2E",X"38",X"10",X"1E",X"00",X"FE",X"F3",X"38",X"36",X"1E",X"E0",X"FE",X"FA",X"38",X"30",
		X"1E",X"EC",X"18",X"2C",X"1E",X"EC",X"FE",X"05",X"38",X"26",X"1E",X"FC",X"FE",X"0A",X"38",X"20",
		X"1E",X"FF",X"FE",X"F3",X"38",X"1A",X"1E",X"1F",X"FE",X"FA",X"38",X"14",X"1E",X"13",X"18",X"10",
		X"1E",X"13",X"FE",X"04",X"38",X"0A",X"1E",X"03",X"FE",X"07",X"38",X"04",X"1E",X"00",X"18",X"00",
		X"21",X"4E",X"5D",X"7A",X"85",X"30",X"01",X"24",X"6F",X"E9",X"7B",X"A2",X"67",X"C9",X"C3",X"72",
		X"5D",X"C3",X"72",X"5D",X"C3",X"AE",X"5D",X"C3",X"E0",X"5D",X"C3",X"10",X"5E",X"C3",X"40",X"5E",
		X"C3",X"40",X"5E",X"C3",X"40",X"5E",X"C3",X"10",X"5E",X"C3",X"E0",X"5D",X"C3",X"AE",X"5D",X"C3",
		X"72",X"5D",X"3A",X"E1",X"F0",X"FE",X"01",X"78",X"28",X"28",X"38",X"10",X"16",X"00",X"FE",X"F1",
		X"38",X"C8",X"16",X"86",X"FE",X"F8",X"38",X"C2",X"16",X"96",X"18",X"BE",X"16",X"9F",X"FE",X"07",
		X"38",X"B8",X"16",X"FF",X"FE",X"F0",X"38",X"B2",X"16",X"79",X"FE",X"F6",X"38",X"AC",X"16",X"69",
		X"18",X"A8",X"16",X"60",X"FE",X"07",X"DA",X"4A",X"5D",X"16",X"00",X"C3",X"4A",X"5D",X"3A",X"E1",
		X"F0",X"FE",X"01",X"28",X"26",X"78",X"38",X"10",X"16",X"00",X"FE",X"F1",X"38",X"8C",X"16",X"86",
		X"FE",X"FB",X"38",X"86",X"16",X"96",X"18",X"82",X"16",X"FF",X"FE",X"F1",X"DA",X"4A",X"5D",X"16",
		X"79",X"FE",X"FB",X"DA",X"4A",X"5D",X"16",X"69",X"C3",X"4A",X"5D",X"16",X"00",X"C3",X"4A",X"5D",
		X"3A",X"E1",X"F0",X"FE",X"01",X"28",X"F4",X"78",X"38",X"13",X"16",X"00",X"FE",X"F1",X"DA",X"4A",
		X"5D",X"16",X"86",X"FE",X"FB",X"DA",X"4A",X"5D",X"16",X"96",X"C3",X"4A",X"5D",X"16",X"FF",X"FE",
		X"F1",X"DA",X"4A",X"5D",X"16",X"39",X"FE",X"FB",X"DA",X"4A",X"5D",X"16",X"09",X"C3",X"4A",X"5D",
		X"3A",X"E1",X"F0",X"FE",X"01",X"28",X"C4",X"78",X"38",X"13",X"16",X"00",X"FE",X"F1",X"DA",X"4A",
		X"5D",X"16",X"E6",X"FE",X"F8",X"DA",X"4A",X"5D",X"16",X"F6",X"C3",X"4A",X"5D",X"16",X"FF",X"FE",
		X"F1",X"DA",X"4A",X"5D",X"16",X"19",X"FE",X"FA",X"DA",X"4A",X"5D",X"16",X"09",X"C3",X"4A",X"5D",
		X"3A",X"E1",X"F0",X"FE",X"01",X"28",X"94",X"78",X"38",X"1A",X"16",X"00",X"FE",X"ED",X"DA",X"4A",
		X"5D",X"16",X"E0",X"FE",X"F2",X"DA",X"4A",X"5D",X"16",X"E6",X"FE",X"FD",X"DA",X"4A",X"5D",X"16",
		X"F6",X"C3",X"4A",X"5D",X"16",X"FF",X"FE",X"EC",X"DA",X"4A",X"5D",X"16",X"1F",X"FE",X"F1",X"DA",
		X"4A",X"5D",X"16",X"19",X"FE",X"FC",X"DA",X"4A",X"5D",X"16",X"09",X"C3",X"4A",X"5D",X"3A",X"E8",
		X"F0",X"FE",X"01",X"30",X"1A",X"3A",X"E7",X"F0",X"FE",X"01",X"D8",X"20",X"03",X"32",X"E8",X"F0",
		X"3D",X"47",X"3A",X"03",X"F0",X"E6",X"03",X"78",X"28",X"01",X"AF",X"32",X"E7",X"F0",X"C9",X"20",
		X"5B",X"3A",X"00",X"F0",X"B7",X"C8",X"D6",X"08",X"47",X"3E",X"0C",X"CB",X"40",X"28",X"02",X"ED",
		X"44",X"80",X"32",X"E2",X"F0",X"AF",X"32",X"E1",X"F0",X"3C",X"32",X"D9",X"F0",X"3C",X"32",X"E8",
		X"F0",X"0E",X"29",X"CD",X"4E",X"3D",X"3A",X"FC",X"F0",X"32",X"FD",X"F0",X"3C",X"32",X"FC",X"F0",
		X"21",X"E4",X"F0",X"36",X"C0",X"21",X"E3",X"F0",X"36",X"01",X"21",X"DB",X"F0",X"36",X"09",X"3A",
		X"82",X"F0",X"C6",X"02",X"32",X"E0",X"F0",X"AF",X"32",X"DF",X"F0",X"32",X"DE",X"F0",X"32",X"E9",
		X"F0",X"32",X"EB",X"F0",X"32",X"EC",X"F0",X"32",X"EA",X"F0",X"18",X"0A",X"3A",X"F3",X"F0",X"B7",
		X"28",X"04",X"3D",X"32",X"F3",X"F0",X"3A",X"E3",X"F0",X"47",X"3A",X"82",X"F0",X"21",X"E0",X"F0",
		X"96",X"4F",X"21",X"E4",X"F0",X"CB",X"7F",X"28",X"06",X"86",X"38",X"10",X"05",X"18",X"04",X"86",
		X"30",X"0A",X"04",X"20",X"07",X"C5",X"0E",X"2B",X"CD",X"4E",X"3D",X"C1",X"77",X"78",X"32",X"E3",
		X"F0",X"B7",X"CA",X"BC",X"5F",X"47",X"3A",X"E8",X"F0",X"FE",X"04",X"CA",X"BC",X"5F",X"3A",X"E9",
		X"F0",X"B7",X"78",X"20",X"37",X"FE",X"FF",X"20",X"73",X"3A",X"E4",X"F0",X"FE",X"80",X"30",X"6C",
		X"3A",X"E8",X"F0",X"FE",X"03",X"28",X"58",X"21",X"E9",X"F0",X"36",X"01",X"21",X"DB",X"F0",X"36",
		X"03",X"3A",X"82",X"F0",X"D6",X"02",X"32",X"E0",X"F0",X"36",X"02",X"AF",X"32",X"DF",X"F0",X"32",
		X"DE",X"F0",X"32",X"EB",X"F0",X"3A",X"00",X"F0",X"32",X"E2",X"F0",X"C9",X"FE",X"01",X"20",X"3C",
		X"3A",X"E4",X"F0",X"FE",X"C0",X"38",X"35",X"3A",X"E8",X"F0",X"FE",X"03",X"28",X"21",X"21",X"DB",
		X"F0",X"36",X"09",X"3A",X"82",X"F0",X"C6",X"02",X"32",X"E0",X"F0",X"AF",X"32",X"DF",X"F0",X"32",
		X"DE",X"F0",X"32",X"E9",X"F0",X"32",X"EB",X"F0",X"3A",X"00",X"F0",X"32",X"E2",X"F0",X"C9",X"AF",
		X"32",X"E8",X"F0",X"32",X"D9",X"F0",X"0E",X"2C",X"CD",X"4E",X"3D",X"C9",X"3A",X"E1",X"F0",X"47",
		X"3A",X"DE",X"F0",X"B7",X"28",X"16",X"21",X"E2",X"F0",X"CB",X"7F",X"28",X"06",X"86",X"38",X"07",
		X"05",X"18",X"04",X"86",X"30",X"01",X"04",X"77",X"78",X"32",X"E1",X"F0",X"3A",X"E8",X"F0",X"FE",
		X"04",X"C8",X"3A",X"03",X"F0",X"E6",X"13",X"28",X"06",X"21",X"E8",X"F0",X"36",X"03",X"C9",X"3A",
		X"E8",X"F0",X"FE",X"03",X"CA",X"FA",X"61",X"3A",X"E9",X"F0",X"B7",X"C2",X"82",X"60",X"3A",X"E3",
		X"F0",X"FE",X"01",X"20",X"29",X"CB",X"79",X"C2",X"E4",X"60",X"3A",X"E4",X"F0",X"FE",X"80",X"38",
		X"0A",X"3A",X"82",X"F0",X"3C",X"32",X"E0",X"F0",X"C3",X"E4",X"60",X"3A",X"DF",X"F0",X"21",X"DD",
		X"F0",X"86",X"30",X"04",X"21",X"E0",X"F0",X"34",X"32",X"DF",X"F0",X"C3",X"E4",X"60",X"30",X"3C",
		X"3A",X"82",X"F0",X"B7",X"20",X"1C",X"3A",X"00",X"F0",X"D6",X"08",X"21",X"E2",X"F0",X"96",X"30",
		X"02",X"ED",X"44",X"FE",X"11",X"30",X"0B",X"FE",X"0A",X"38",X"07",X"3A",X"E4",X"F0",X"FE",X"E8",
		X"38",X"1A",X"21",X"E4",X"F0",X"3A",X"01",X"F0",X"D6",X"20",X"96",X"38",X"A8",X"7E",X"FE",X"40",
		X"30",X"0A",X"3A",X"EB",X"F0",X"B7",X"20",X"04",X"3C",X"32",X"EB",X"F0",X"CB",X"79",X"28",X"74",
		X"3A",X"DF",X"F0",X"21",X"DD",X"F0",X"96",X"30",X"04",X"21",X"E0",X"F0",X"35",X"32",X"DF",X"F0",
		X"18",X"62",X"3A",X"E3",X"F0",X"FE",X"01",X"20",X"21",X"3A",X"EB",X"F0",X"B7",X"20",X"04",X"3C",
		X"32",X"EB",X"F0",X"79",X"CB",X"7F",X"28",X"38",X"3A",X"DF",X"F0",X"21",X"DD",X"F0",X"96",X"30",
		X"04",X"21",X"E0",X"F0",X"35",X"32",X"DF",X"F0",X"18",X"3A",X"30",X"0B",X"21",X"E4",X"F0",X"3A",
		X"01",X"F0",X"C6",X"28",X"96",X"38",X"D2",X"79",X"D6",X"02",X"CB",X"7F",X"28",X"12",X"3A",X"DF",
		X"F0",X"21",X"DD",X"F0",X"96",X"30",X"04",X"21",X"E0",X"F0",X"35",X"32",X"DF",X"F0",X"18",X"14",
		X"FE",X"03",X"38",X"10",X"3A",X"DF",X"F0",X"21",X"DD",X"F0",X"86",X"30",X"04",X"21",X"E0",X"F0",
		X"34",X"32",X"DF",X"F0",X"3A",X"EB",X"F0",X"B7",X"C2",X"2C",X"62",X"3A",X"00",X"F0",X"D6",X"08",
		X"47",X"3A",X"E3",X"F0",X"B7",X"20",X"61",X"3A",X"E1",X"F0",X"B7",X"20",X"5B",X"21",X"E4",X"F0",
		X"3A",X"82",X"F0",X"B7",X"3A",X"01",X"F0",X"20",X"02",X"C6",X"14",X"96",X"38",X"4A",X"7E",X"FE",
		X"20",X"38",X"45",X"78",X"21",X"E2",X"F0",X"96",X"30",X"02",X"ED",X"44",X"FE",X"11",X"30",X"38",
		X"FE",X"0A",X"38",X"34",X"3A",X"19",X"F0",X"21",X"18",X"F0",X"B6",X"20",X"2B",X"3A",X"EE",X"F0",
		X"21",X"EF",X"F0",X"B6",X"20",X"22",X"3A",X"F3",X"F0",X"B7",X"20",X"1C",X"3A",X"FD",X"F0",X"B7",
		X"28",X"16",X"3D",X"32",X"FD",X"F0",X"21",X"EE",X"F0",X"36",X"01",X"21",X"F3",X"F0",X"36",X"30",
		X"20",X"06",X"21",X"E8",X"F0",X"36",X"03",X"C9",X"21",X"EA",X"F0",X"7E",X"B7",X"28",X"02",X"35",
		X"C9",X"36",X"0C",X"3A",X"E9",X"F0",X"B7",X"20",X"3C",X"16",X"FF",X"1E",X"08",X"3A",X"E1",X"F0",
		X"FE",X"01",X"38",X"08",X"28",X"5F",X"16",X"01",X"1E",X"0A",X"18",X"59",X"3A",X"E2",X"F0",X"0E",
		X"0A",X"90",X"30",X"08",X"ED",X"44",X"0E",X"08",X"16",X"01",X"1E",X"0A",X"FE",X"11",X"30",X"45",
		X"FE",X"0A",X"30",X"07",X"7A",X"ED",X"44",X"57",X"59",X"18",X"3A",X"AF",X"32",X"DE",X"F0",X"3E",
		X"09",X"32",X"DB",X"F0",X"C9",X"16",X"FF",X"1E",X"04",X"3A",X"E1",X"F0",X"FE",X"01",X"38",X"08",
		X"28",X"23",X"16",X"01",X"1E",X"02",X"18",X"1D",X"3A",X"E2",X"F0",X"0E",X"02",X"90",X"30",X"08",
		X"ED",X"44",X"0E",X"04",X"16",X"01",X"1E",X"02",X"FE",X"11",X"30",X"09",X"FE",X"0A",X"30",X"20",
		X"7A",X"ED",X"44",X"57",X"59",X"21",X"DB",X"F0",X"7B",X"BE",X"C8",X"7A",X"32",X"DE",X"F0",X"16",
		X"03",X"3A",X"E9",X"F0",X"B7",X"20",X"02",X"16",X"09",X"7E",X"BA",X"28",X"01",X"5A",X"73",X"C9",
		X"AF",X"32",X"DE",X"F0",X"3E",X"03",X"32",X"DB",X"F0",X"C9",X"3A",X"E9",X"F0",X"B7",X"20",X"15",
		X"0C",X"CB",X"79",X"C0",X"3A",X"DF",X"F0",X"21",X"DD",X"F0",X"86",X"30",X"04",X"21",X"E0",X"F0",
		X"34",X"32",X"DF",X"F0",X"C9",X"79",X"D6",X"02",X"CB",X"7F",X"C8",X"3A",X"DF",X"F0",X"21",X"DD",
		X"F0",X"96",X"30",X"04",X"21",X"E0",X"F0",X"35",X"32",X"DF",X"F0",X"C9",X"47",X"3A",X"EC",X"F0",
		X"B7",X"28",X"05",X"3D",X"32",X"EC",X"F0",X"C9",X"78",X"FE",X"01",X"20",X"34",X"3A",X"E9",X"F0",
		X"B7",X"20",X"16",X"3A",X"E2",X"F0",X"FE",X"80",X"38",X"08",X"3E",X"0C",X"21",X"DB",X"F0",X"96",
		X"18",X"1B",X"3A",X"DB",X"F0",X"C6",X"02",X"18",X"14",X"3A",X"E2",X"F0",X"FE",X"80",X"38",X"07",
		X"3A",X"DB",X"F0",X"C6",X"10",X"18",X"06",X"3E",X"1E",X"21",X"DB",X"F0",X"96",X"32",X"EB",X"F0",
		X"C9",X"D6",X"02",X"CB",X"27",X"CB",X"27",X"21",X"9E",X"62",X"85",X"30",X"01",X"24",X"6F",X"7E",
		X"32",X"DB",X"F0",X"23",X"7E",X"32",X"DE",X"F0",X"23",X"7E",X"32",X"EC",X"F0",X"23",X"7E",X"32",
		X"EB",X"F0",X"B7",X"C0",X"3A",X"E9",X"F0",X"2F",X"E6",X"01",X"32",X"E9",X"F0",X"C9",X"09",X"01",
		X"08",X"03",X"08",X"00",X"08",X"04",X"07",X"FF",X"08",X"05",X"06",X"FE",X"08",X"06",X"05",X"FD",
		X"08",X"07",X"04",X"FE",X"08",X"08",X"03",X"FF",X"08",X"09",X"03",X"00",X"08",X"00",X"09",X"FF",
		X"08",X"0B",X"0A",X"00",X"08",X"0C",X"0B",X"01",X"08",X"0D",X"00",X"02",X"08",X"0E",X"01",X"03",
		X"08",X"0F",X"02",X"02",X"08",X"10",X"03",X"01",X"08",X"11",X"03",X"00",X"08",X"00",X"03",X"01",
		X"08",X"13",X"04",X"00",X"08",X"14",X"05",X"FF",X"08",X"15",X"06",X"FE",X"08",X"16",X"07",X"FD",
		X"08",X"17",X"08",X"FE",X"08",X"18",X"09",X"FF",X"08",X"19",X"09",X"00",X"08",X"00",X"03",X"FF",
		X"08",X"1B",X"02",X"00",X"08",X"1C",X"01",X"01",X"08",X"1D",X"00",X"02",X"08",X"1E",X"0B",X"03",
		X"08",X"1F",X"0A",X"02",X"08",X"20",X"09",X"01",X"08",X"21",X"09",X"00",X"08",X"00",X"3A",X"EE",
		X"F0",X"B7",X"C8",X"FD",X"21",X"D8",X"F9",X"3D",X"47",X"CB",X"27",X"80",X"21",X"3D",X"63",X"85",
		X"30",X"01",X"24",X"6F",X"E9",X"AF",X"FD",X"77",X"00",X"32",X"EE",X"F0",X"C9",X"C3",X"46",X"63",
		X"C3",X"6F",X"63",X"C3",X"BC",X"63",X"3A",X"E3",X"F0",X"B7",X"20",X"E9",X"3A",X"00",X"F0",X"21",
		X"E2",X"F0",X"96",X"0E",X"01",X"30",X"04",X"0E",X"00",X"ED",X"44",X"FE",X"28",X"D2",X"35",X"63",
		X"21",X"EE",X"F0",X"36",X"02",X"21",X"F0",X"F0",X"36",X"08",X"21",X"F2",X"F0",X"71",X"C9",X"3A",
		X"E3",X"F0",X"B7",X"20",X"C0",X"21",X"F0",X"F0",X"35",X"28",X"29",X"3A",X"F2",X"F0",X"B7",X"3A",
		X"E2",X"F0",X"20",X"0A",X"3C",X"FD",X"77",X"00",X"FD",X"36",X"01",X"20",X"18",X"09",X"C6",X"10",
		X"FD",X"77",X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"01",X"3A",X"E4",X"F0",X"C6",X"F5",
		X"FD",X"77",X"03",X"C9",X"36",X"02",X"3A",X"00",X"F0",X"21",X"E2",X"F0",X"96",X"30",X"02",X"ED",
		X"44",X"FE",X"30",X"D2",X"35",X"63",X"21",X"EE",X"F0",X"36",X"03",X"C9",X"3A",X"E3",X"F0",X"B7",
		X"C2",X"35",X"63",X"21",X"F0",X"F0",X"35",X"28",X"29",X"3A",X"F2",X"F0",X"B7",X"3A",X"E2",X"F0",
		X"20",X"0A",X"3C",X"FD",X"77",X"00",X"FD",X"36",X"01",X"20",X"18",X"09",X"C6",X"10",X"FD",X"77",
		X"00",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"02",X"3A",X"E4",X"F0",X"C6",X"F5",X"FD",X"77",
		X"03",X"C9",X"36",X"18",X"3A",X"F2",X"F0",X"B7",X"3A",X"E2",X"F0",X"20",X"04",X"C6",X"F8",X"18",
		X"02",X"C6",X"1A",X"32",X"F4",X"F0",X"DD",X"21",X"C0",X"F9",X"DD",X"77",X"00",X"3A",X"E4",X"F0",
		X"C6",X"F9",X"32",X"F5",X"F0",X"DD",X"77",X"03",X"DD",X"36",X"02",X"68",X"AF",X"32",X"F6",X"F0",
		X"32",X"EE",X"F0",X"FD",X"77",X"00",X"3C",X"32",X"EF",X"F0",X"3A",X"DE",X"F0",X"B7",X"28",X"08",
		X"CB",X"7F",X"28",X"03",X"3C",X"18",X"01",X"3D",X"32",X"F7",X"F0",X"3A",X"E0",X"F0",X"B7",X"28",
		X"08",X"CB",X"7F",X"28",X"03",X"3C",X"18",X"01",X"3D",X"32",X"F8",X"F0",X"0E",X"0D",X"CD",X"4E",
		X"3D",X"C9",X"3A",X"51",X"F0",X"B7",X"C8",X"16",X"06",X"DD",X"21",X"8B",X"F2",X"DD",X"7E",X"01",
		X"47",X"E6",X"40",X"CA",X"C9",X"66",X"78",X"E6",X"0A",X"C2",X"7F",X"66",X"78",X"E6",X"04",X"28",
		X"08",X"DD",X"7E",X"0C",X"FE",X"70",X"D2",X"7F",X"66",X"DD",X"7E",X"07",X"FE",X"D0",X"D2",X"7F",
		X"66",X"FE",X"30",X"DA",X"7F",X"66",X"26",X"F4",X"2E",X"F4",X"DD",X"7E",X"13",X"B7",X"28",X"21",
		X"26",X"03",X"47",X"DD",X"4E",X"12",X"C5",X"FD",X"E1",X"DD",X"7E",X"05",X"D6",X"0B",X"FD",X"77",
		X"00",X"FD",X"7E",X"01",X"EE",X"10",X"FD",X"77",X"01",X"DD",X"7E",X"07",X"C6",X"02",X"FD",X"77",
		X"03",X"DD",X"7E",X"15",X"B7",X"28",X"21",X"2E",X"03",X"47",X"DD",X"4E",X"14",X"C5",X"FD",X"E1",
		X"DD",X"7E",X"05",X"C6",X"0C",X"FD",X"77",X"00",X"FD",X"7E",X"01",X"EE",X"10",X"FD",X"77",X"01",
		X"DD",X"7E",X"07",X"C6",X"02",X"FD",X"77",X"03",X"3A",X"03",X"F0",X"E6",X"10",X"C2",X"95",X"65",
		X"3A",X"01",X"F0",X"47",X"3A",X"04",X"F0",X"80",X"D6",X"0C",X"DD",X"BE",X"07",X"DA",X"95",X"65",
		X"DD",X"7E",X"07",X"DD",X"86",X"0E",X"D6",X"0C",X"B8",X"DA",X"95",X"65",X"3A",X"00",X"F0",X"47",
		X"C6",X"10",X"84",X"DD",X"BE",X"05",X"DA",X"95",X"65",X"DD",X"7E",X"05",X"B8",X"30",X"33",X"C6",
		X"10",X"85",X"B8",X"DA",X"95",X"65",X"DD",X"7E",X"15",X"B7",X"CA",X"C9",X"66",X"67",X"DD",X"6E",
		X"14",X"36",X"00",X"DD",X"36",X"15",X"00",X"DD",X"7E",X"13",X"B7",X"20",X"3F",X"DD",X"7E",X"01",
		X"EE",X"40",X"DD",X"77",X"01",X"21",X"51",X"F0",X"35",X"20",X"31",X"0E",X"32",X"CD",X"4E",X"3D",
		X"18",X"2A",X"DD",X"7E",X"13",X"B7",X"CA",X"C9",X"66",X"67",X"DD",X"6E",X"12",X"36",X"00",X"DD",
		X"36",X"13",X"00",X"DD",X"7E",X"15",X"B7",X"20",X"13",X"DD",X"7E",X"01",X"EE",X"40",X"DD",X"77",
		X"01",X"21",X"51",X"F0",X"35",X"20",X"05",X"0E",X"32",X"CD",X"4E",X"3D",X"3A",X"03",X"F0",X"F6",
		X"02",X"32",X"03",X"F0",X"3A",X"00",X"F0",X"DD",X"BE",X"05",X"3E",X"02",X"06",X"07",X"30",X"04",
		X"ED",X"44",X"06",X"00",X"32",X"A1",X"F0",X"21",X"02",X"F0",X"70",X"0E",X"35",X"CD",X"4E",X"3D",
		X"DD",X"36",X"04",X"00",X"C9",X"1E",X"06",X"FD",X"21",X"8B",X"F2",X"FD",X"7E",X"00",X"DD",X"BE",
		X"00",X"CA",X"74",X"66",X"FD",X"7E",X"01",X"E6",X"80",X"CA",X"74",X"66",X"FD",X"7E",X"08",X"B7",
		X"C2",X"74",X"66",X"FD",X"7E",X"07",X"47",X"FD",X"86",X"0E",X"D6",X"04",X"DD",X"BE",X"07",X"DA",
		X"74",X"66",X"DD",X"7E",X"07",X"DD",X"86",X"0E",X"D6",X"04",X"B8",X"DA",X"74",X"66",X"FD",X"7E",
		X"05",X"47",X"C6",X"10",X"84",X"DD",X"BE",X"05",X"DA",X"74",X"66",X"DD",X"7E",X"05",X"B8",X"30",
		X"33",X"C6",X"10",X"85",X"B8",X"DA",X"74",X"66",X"DD",X"7E",X"15",X"B7",X"CA",X"74",X"66",X"67",
		X"DD",X"6E",X"14",X"36",X"00",X"DD",X"36",X"15",X"00",X"DD",X"7E",X"13",X"B7",X"20",X"3E",X"DD",
		X"7E",X"01",X"EE",X"40",X"DD",X"77",X"01",X"21",X"51",X"F0",X"35",X"20",X"30",X"0E",X"32",X"CD",
		X"4E",X"3D",X"18",X"29",X"DD",X"7E",X"13",X"B7",X"28",X"5A",X"67",X"DD",X"6E",X"12",X"36",X"00",
		X"DD",X"36",X"13",X"00",X"DD",X"7E",X"15",X"B7",X"20",X"13",X"DD",X"7E",X"01",X"EE",X"40",X"DD",
		X"77",X"01",X"21",X"51",X"F0",X"35",X"20",X"05",X"0E",X"32",X"CD",X"4E",X"3D",X"FD",X"7E",X"01",
		X"47",X"E6",X"0A",X"C2",X"C9",X"66",X"78",X"E6",X"40",X"20",X"7E",X"FD",X"7E",X"02",X"E6",X"0F",
		X"FE",X"05",X"30",X"75",X"78",X"F6",X"08",X"FD",X"77",X"01",X"FD",X"7E",X"18",X"B7",X"28",X"0A",
		X"67",X"FD",X"6E",X"17",X"36",X"00",X"FD",X"36",X"18",X"00",X"FD",X"36",X"16",X"7F",X"FD",X"36",
		X"0C",X"01",X"18",X"55",X"01",X"23",X"00",X"FD",X"09",X"1D",X"C2",X"9B",X"65",X"18",X"4A",X"DD",
		X"7E",X"01",X"E6",X"40",X"C8",X"DD",X"7E",X"01",X"EE",X"40",X"DD",X"77",X"01",X"DD",X"7E",X"13",
		X"B7",X"28",X"12",X"67",X"DD",X"6E",X"12",X"36",X"00",X"DD",X"36",X"13",X"00",X"DD",X"7E",X"02",
		X"F6",X"20",X"DD",X"77",X"02",X"DD",X"7E",X"15",X"B7",X"28",X"12",X"67",X"DD",X"6E",X"14",X"36",
		X"00",X"DD",X"36",X"15",X"00",X"DD",X"7E",X"02",X"F6",X"40",X"DD",X"77",X"02",X"21",X"51",X"F0",
		X"35",X"20",X"06",X"0E",X"32",X"CD",X"4E",X"3D",X"C9",X"01",X"23",X"00",X"DD",X"09",X"15",X"C2",
		X"5D",X"64",X"C9",X"21",X"B0",X"F0",X"7E",X"E5",X"47",X"CB",X"27",X"80",X"21",X"E5",X"66",X"85",
		X"30",X"01",X"24",X"6F",X"E9",X"C3",X"09",X"67",X"C3",X"F1",X"67",X"C3",X"ED",X"6D",X"C3",X"8E",
		X"6F",X"C3",X"84",X"70",X"C3",X"E2",X"70",X"C3",X"F0",X"70",X"C3",X"1A",X"71",X"C3",X"4B",X"71",
		X"C3",X"AD",X"71",X"C3",X"D9",X"71",X"C3",X"12",X"72",X"AF",X"32",X"28",X"F0",X"32",X"26",X"F0",
		X"3A",X"15",X"F0",X"B7",X"C2",X"D6",X"67",X"3A",X"56",X"F0",X"D6",X"8E",X"20",X"09",X"32",X"07",
		X"F0",X"E1",X"34",X"23",X"36",X"30",X"C9",X"06",X"00",X"0E",X"D0",X"FD",X"21",X"5B",X"F2",X"CD",
		X"B5",X"41",X"3A",X"AF",X"F0",X"B7",X"28",X"0B",X"FD",X"7E",X"02",X"B7",X"28",X"05",X"FD",X"7E",
		X"03",X"18",X"0A",X"FD",X"7E",X"01",X"FE",X"60",X"30",X"03",X"FD",X"7E",X"03",X"C6",X"03",X"32",
		X"07",X"F0",X"FD",X"2A",X"2A",X"F0",X"E1",X"34",X"23",X"3A",X"A1",X"F0",X"B7",X"20",X"18",X"FD",
		X"36",X"02",X"20",X"FD",X"2A",X"2C",X"F0",X"FD",X"36",X"00",X"00",X"36",X"28",X"0E",X"13",X"CD",
		X"4E",X"3D",X"21",X"AD",X"F0",X"35",X"C9",X"3A",X"56",X"F0",X"E6",X"80",X"20",X"08",X"36",X"28",
		X"0E",X"26",X"CD",X"4E",X"3D",X"C9",X"36",X"30",X"FD",X"4E",X"00",X"FD",X"7E",X"03",X"C6",X"0A",
		X"47",X"CD",X"21",X"72",X"06",X"04",X"2B",X"7E",X"FE",X"F0",X"28",X"18",X"FE",X"B0",X"28",X"18",
		X"FE",X"A9",X"28",X"1F",X"FE",X"E9",X"28",X"1B",X"FE",X"E2",X"28",X"1B",X"FE",X"A2",X"28",X"17",
		X"23",X"10",X"E4",X"C9",X"36",X"D5",X"18",X"02",X"36",X"95",X"22",X"9B",X"F0",X"0E",X"13",X"CD",
		X"4E",X"3D",X"C9",X"36",X"E8",X"18",X"02",X"36",X"9F",X"0E",X"13",X"CD",X"4E",X"3D",X"AF",X"32",
		X"56",X"F0",X"32",X"9C",X"F0",X"C9",X"32",X"07",X"F0",X"E1",X"34",X"23",X"36",X"28",X"3A",X"A1",
		X"F0",X"B7",X"C0",X"FD",X"2A",X"2A",X"F0",X"FD",X"36",X"02",X"B7",X"0E",X"13",X"CD",X"4E",X"3D",
		X"C9",X"3A",X"15",X"F0",X"B7",X"C2",X"FC",X"69",X"E1",X"23",X"35",X"7E",X"FE",X"1F",X"DA",X"74",
		X"69",X"FD",X"2A",X"2A",X"F0",X"C2",X"0D",X"69",X"CD",X"70",X"72",X"3A",X"56",X"F0",X"FE",X"8E",
		X"28",X"69",X"E6",X"80",X"20",X"26",X"0E",X"13",X"CD",X"4E",X"3D",X"FD",X"7E",X"00",X"B7",X"C8",
		X"FD",X"7E",X"02",X"FE",X"20",X"C8",X"FD",X"36",X"02",X"20",X"FD",X"2A",X"2C",X"F0",X"FD",X"7E",
		X"00",X"B7",X"C8",X"FD",X"36",X"00",X"00",X"21",X"AD",X"F0",X"35",X"C9",X"FD",X"7E",X"00",X"B7",
		X"20",X"0B",X"3A",X"56",X"F0",X"FE",X"85",X"CA",X"07",X"69",X"3A",X"08",X"F0",X"06",X"F8",X"FE",
		X"F8",X"30",X"28",X"06",X"08",X"FE",X"18",X"38",X"22",X"4F",X"FD",X"7E",X"03",X"C6",X"0A",X"47",
		X"CD",X"21",X"72",X"3A",X"A1",X"F0",X"CB",X"7F",X"06",X"F0",X"28",X"02",X"06",X"B0",X"23",X"7E",
		X"FE",X"AF",X"28",X"07",X"FE",X"EF",X"28",X"03",X"B8",X"20",X"9B",X"21",X"26",X"F0",X"36",X"01",
		X"FD",X"4E",X"03",X"FD",X"7E",X"00",X"B7",X"28",X"15",X"47",X"FD",X"36",X"00",X"00",X"FD",X"2A",
		X"2C",X"F0",X"FD",X"36",X"00",X"00",X"3A",X"AD",X"F0",X"D6",X"02",X"32",X"AD",X"F0",X"11",X"04",
		X"00",X"FD",X"21",X"78",X"F8",X"FD",X"36",X"02",X"64",X"FD",X"36",X"01",X"00",X"79",X"D6",X"10",
		X"FD",X"77",X"03",X"78",X"C6",X"08",X"FD",X"77",X"00",X"FD",X"19",X"FD",X"77",X"00",X"FD",X"36",
		X"02",X"65",X"FD",X"36",X"01",X"00",X"FD",X"71",X"03",X"FD",X"19",X"FD",X"36",X"02",X"66",X"FD",
		X"36",X"01",X"00",X"79",X"D6",X"10",X"FD",X"77",X"03",X"78",X"D6",X"08",X"FD",X"77",X"00",X"FD",
		X"19",X"FD",X"77",X"00",X"FD",X"36",X"02",X"67",X"FD",X"36",X"01",X"00",X"FD",X"71",X"03",X"FD",
		X"19",X"FD",X"70",X"00",X"FD",X"36",X"02",X"5E",X"FD",X"36",X"01",X"00",X"79",X"D6",X"06",X"FD",
		X"77",X"03",X"0E",X"14",X"CD",X"4E",X"3D",X"0E",X"33",X"CD",X"4E",X"3D",X"C9",X"FE",X"2A",X"20",
		X"14",X"3A",X"9C",X"F0",X"B7",X"28",X"0E",X"2A",X"9B",X"F0",X"7E",X"FE",X"D5",X"28",X"04",X"FE",
		X"95",X"20",X"02",X"36",X"EF",X"FD",X"7E",X"03",X"D6",X"03",X"38",X"2B",X"FD",X"77",X"03",X"3A",
		X"A1",X"F0",X"FD",X"86",X"00",X"FE",X"05",X"38",X"21",X"FE",X"FB",X"30",X"1D",X"FD",X"77",X"00",
		X"47",X"FD",X"7E",X"02",X"FE",X"20",X"C8",X"FD",X"2A",X"2C",X"F0",X"FD",X"70",X"00",X"FD",X"7E",
		X"03",X"D6",X"03",X"FD",X"77",X"03",X"C9",X"FD",X"7E",X"00",X"32",X"08",X"F0",X"FD",X"36",X"00",
		X"00",X"FD",X"2A",X"2C",X"F0",X"FD",X"36",X"00",X"00",X"36",X"20",X"3A",X"AD",X"F0",X"D6",X"02",
		X"32",X"AD",X"F0",X"C9",X"B7",X"20",X"0D",X"2B",X"34",X"0E",X"14",X"CD",X"4E",X"3D",X"21",X"25",
		X"F0",X"36",X"00",X"C9",X"47",X"3A",X"26",X"F0",X"B7",X"28",X"65",X"78",X"FE",X"16",X"20",X"34",
		X"11",X"04",X"00",X"FD",X"21",X"78",X"F8",X"FD",X"36",X"00",X"00",X"FD",X"36",X"03",X"00",X"FD",
		X"19",X"FD",X"36",X"00",X"00",X"FD",X"36",X"03",X"00",X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",
		X"36",X"03",X"00",X"FD",X"19",X"FD",X"36",X"00",X"00",X"FD",X"36",X"03",X"00",X"FD",X"19",X"FD",
		X"36",X"02",X"5F",X"C9",X"FE",X"0F",X"20",X"09",X"FD",X"21",X"88",X"F8",X"FD",X"36",X"02",X"60",
		X"C9",X"FE",X"08",X"20",X"09",X"FD",X"21",X"88",X"F8",X"FD",X"36",X"02",X"61",X"C9",X"FE",X"01",
		X"C0",X"AF",X"FD",X"21",X"88",X"F8",X"FD",X"77",X"00",X"FD",X"77",X"03",X"32",X"26",X"F0",X"C9",
		X"FD",X"2A",X"2A",X"F0",X"FD",X"7E",X"00",X"B7",X"C8",X"C3",X"39",X"6B",X"E1",X"23",X"35",X"7E",
		X"FE",X"1F",X"DA",X"19",X"6B",X"CA",X"0F",X"6A",X"FD",X"2A",X"2A",X"F0",X"C3",X"25",X"69",X"DD",
		X"2A",X"2A",X"F0",X"DD",X"7E",X"00",X"B7",X"28",X"5F",X"CD",X"70",X"72",X"3A",X"0A",X"F0",X"B7",
		X"28",X"07",X"3A",X"56",X"F0",X"E6",X"01",X"18",X"35",X"3A",X"56",X"F0",X"FE",X"01",X"28",X"04",
		X"FE",X"09",X"20",X"04",X"3E",X"01",X"18",X"26",X"06",X"00",X"DD",X"4E",X"03",X"FD",X"21",X"5B",
		X"F2",X"CD",X"B5",X"41",X"DD",X"46",X"00",X"CD",X"62",X"45",X"47",X"3E",X"01",X"38",X"0F",X"16",
		X"02",X"79",X"B7",X"20",X"02",X"14",X"78",X"FE",X"0C",X"3E",X"00",X"30",X"01",X"82",X"32",X"26",
		X"F0",X"B7",X"20",X"1A",X"DD",X"36",X"02",X"BF",X"DD",X"2A",X"2C",X"F0",X"DD",X"36",X"02",X"C0",
		X"DD",X"7E",X"03",X"D6",X"04",X"DD",X"77",X"03",X"0E",X"13",X"CD",X"4E",X"3D",X"C9",X"DD",X"36",
		X"02",X"B7",X"FE",X"02",X"20",X"0C",X"DD",X"36",X"01",X"20",X"DD",X"2A",X"2C",X"F0",X"DD",X"36",
		X"01",X"20",X"FD",X"21",X"48",X"F8",X"11",X"04",X"00",X"DD",X"7E",X"00",X"C6",X"08",X"FD",X"77",
		X"00",X"47",X"DD",X"7E",X"03",X"D6",X"04",X"FD",X"77",X"03",X"4F",X"FD",X"36",X"02",X"64",X"FD",
		X"36",X"01",X"00",X"FD",X"19",X"FD",X"70",X"00",X"C6",X"10",X"FD",X"77",X"03",X"FD",X"36",X"02",
		X"65",X"FD",X"36",X"01",X"00",X"FD",X"19",X"78",X"D6",X"10",X"FD",X"77",X"00",X"FD",X"71",X"03",
		X"FD",X"36",X"02",X"64",X"FD",X"36",X"01",X"20",X"FD",X"19",X"FD",X"77",X"00",X"79",X"C6",X"10",
		X"FD",X"77",X"03",X"FD",X"36",X"02",X"65",X"FD",X"36",X"01",X"20",X"FD",X"19",X"DD",X"46",X"00",
		X"FD",X"70",X"00",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"FD",X"36",X"02",X"B7",X"FD",X"36",X"01",
		X"00",X"FD",X"19",X"FD",X"70",X"00",X"C6",X"10",X"FD",X"77",X"03",X"FD",X"36",X"02",X"85",X"FD",
		X"36",X"01",X"00",X"0E",X"33",X"CD",X"4E",X"3D",X"C9",X"B7",X"20",X"0C",X"2B",X"34",X"0E",X"14",
		X"CD",X"4E",X"3D",X"AF",X"32",X"25",X"F0",X"C9",X"FD",X"2A",X"2A",X"F0",X"47",X"FD",X"7E",X"00",
		X"B7",X"C8",X"3A",X"26",X"F0",X"B7",X"C2",X"70",X"6D",X"DD",X"21",X"78",X"F8",X"11",X"04",X"00",
		X"3E",X"1E",X"90",X"47",X"CB",X"27",X"80",X"21",X"5D",X"6B",X"85",X"30",X"01",X"24",X"6F",X"01",
		X"00",X"00",X"3A",X"15",X"F0",X"B7",X"20",X"04",X"06",X"04",X"0E",X"F4",X"E9",X"C3",X"B7",X"6B",
		X"C3",X"B7",X"6B",X"C3",X"D2",X"6B",X"C3",X"D2",X"6B",X"C3",X"D2",X"6B",X"C3",X"F5",X"6B",X"C3",
		X"F5",X"6B",X"C3",X"F5",X"6B",X"C3",X"23",X"6C",X"C3",X"23",X"6C",X"C3",X"23",X"6C",X"C3",X"37",
		X"6C",X"C3",X"37",X"6C",X"C3",X"37",X"6C",X"C3",X"55",X"6C",X"C3",X"55",X"6C",X"C3",X"55",X"6C",
		X"C3",X"82",X"6C",X"C3",X"82",X"6C",X"C3",X"82",X"6C",X"C3",X"AB",X"6C",X"C3",X"AB",X"6C",X"C3",
		X"AB",X"6C",X"C3",X"FA",X"6C",X"C3",X"FA",X"6C",X"C3",X"FA",X"6C",X"C3",X"2F",X"6D",X"C3",X"2F",
		X"6D",X"C3",X"2F",X"6D",X"C3",X"50",X"6D",X"FD",X"7E",X"00",X"80",X"D6",X"04",X"DD",X"77",X"00",
		X"FD",X"7E",X"03",X"81",X"C6",X"08",X"DD",X"77",X"03",X"DD",X"36",X"02",X"35",X"DD",X"36",X"01",
		X"00",X"C9",X"FD",X"7E",X"00",X"80",X"D6",X"04",X"DD",X"77",X"00",X"FD",X"7E",X"03",X"81",X"C6",
		X"04",X"DD",X"77",X"03",X"DD",X"36",X"02",X"36",X"DD",X"36",X"04",X"00",X"DD",X"36",X"06",X"37",
		X"DD",X"36",X"05",X"00",X"C9",X"FD",X"7E",X"00",X"80",X"D6",X"02",X"DD",X"77",X"00",X"47",X"FD",
		X"7E",X"03",X"81",X"DD",X"77",X"03",X"4F",X"DD",X"7E",X"01",X"EE",X"20",X"DD",X"77",X"01",X"DD",
		X"19",X"DD",X"70",X"00",X"79",X"C6",X"0C",X"DD",X"77",X"03",X"DD",X"7E",X"01",X"EE",X"20",X"DD",
		X"77",X"01",X"C9",X"CD",X"F5",X"6B",X"DD",X"19",X"DD",X"70",X"00",X"DD",X"71",X"03",X"DD",X"36",
		X"02",X"18",X"DD",X"36",X"01",X"10",X"C9",X"CD",X"23",X"6C",X"DD",X"36",X"01",X"30",X"DD",X"19",
		X"78",X"D6",X"02",X"DD",X"77",X"00",X"79",X"D6",X"07",X"DD",X"77",X"03",X"DD",X"36",X"02",X"19",
		X"DD",X"36",X"01",X"20",X"C9",X"CD",X"23",X"6C",X"DD",X"36",X"01",X"10",X"DD",X"19",X"78",X"D6",
		X"04",X"DD",X"77",X"00",X"79",X"D6",X"07",X"DD",X"77",X"03",X"DD",X"36",X"01",X"00",X"DD",X"19",
		X"DD",X"77",X"03",X"78",X"C6",X"04",X"DD",X"77",X"00",X"DD",X"36",X"02",X"19",X"DD",X"36",X"01",
		X"10",X"C9",X"CD",X"23",X"6C",X"DD",X"36",X"01",X"30",X"DD",X"19",X"78",X"D6",X"05",X"DD",X"77",
		X"00",X"79",X"D6",X"0B",X"DD",X"77",X"03",X"DD",X"36",X"01",X"30",X"DD",X"19",X"DD",X"77",X"03",
		X"78",X"C6",X"05",X"DD",X"77",X"00",X"DD",X"36",X"01",X"20",X"C9",X"DD",X"36",X"00",X"00",X"DD",
		X"19",X"FD",X"7E",X"00",X"80",X"D6",X"02",X"47",X"DD",X"77",X"00",X"FD",X"7E",X"03",X"81",X"4F",
		X"C6",X"0C",X"DD",X"77",X"03",X"DD",X"36",X"02",X"36",X"DD",X"19",X"DD",X"70",X"00",X"79",X"D6",
		X"04",X"DD",X"77",X"03",X"DD",X"36",X"01",X"10",X"DD",X"19",X"78",X"D6",X"05",X"DD",X"77",X"00",
		X"79",X"D6",X"0B",X"DD",X"77",X"03",X"DD",X"36",X"01",X"20",X"DD",X"19",X"DD",X"77",X"03",X"78",
		X"C6",X"05",X"DD",X"77",X"00",X"DD",X"36",X"01",X"10",X"C9",X"DD",X"19",X"DD",X"36",X"00",X"00",
		X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",X"19",X"FD",X"7E",X"00",X"80",X"47",X"D6",X"07",X"DD",
		X"77",X"00",X"FD",X"7E",X"03",X"81",X"D6",X"0D",X"DD",X"77",X"03",X"DD",X"36",X"01",X"10",X"DD",
		X"19",X"DD",X"77",X"03",X"78",X"C6",X"03",X"DD",X"77",X"00",X"DD",X"36",X"01",X"30",X"C9",X"DD",
		X"21",X"84",X"F8",X"DD",X"36",X"00",X"00",X"DD",X"19",X"FD",X"7E",X"00",X"80",X"D6",X"05",X"DD",
		X"77",X"00",X"FD",X"7E",X"03",X"81",X"D6",X"0D",X"DD",X"77",X"03",X"DD",X"36",X"01",X"10",X"C9",
		X"DD",X"21",X"88",X"F8",X"DD",X"36",X"00",X"00",X"3A",X"15",X"F0",X"B7",X"C0",X"3A",X"56",X"F0",
		X"E6",X"80",X"C8",X"FD",X"2A",X"2A",X"F0",X"FD",X"36",X"00",X"00",X"21",X"AD",X"F0",X"35",X"C9",
		X"78",X"DD",X"2A",X"2C",X"F0",X"FE",X"19",X"20",X"32",X"DD",X"36",X"02",X"B8",X"FD",X"36",X"02",
		X"B7",X"DD",X"21",X"48",X"F8",X"11",X"04",X"00",X"DD",X"36",X"00",X"00",X"DD",X"19",X"DD",X"36",
		X"00",X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",X"19",
		X"DD",X"36",X"00",X"00",X"DD",X"19",X"DD",X"36",X"00",X"00",X"C9",X"FE",X"13",X"20",X"09",X"FD",
		X"36",X"02",X"B9",X"DD",X"36",X"02",X"BA",X"C9",X"FE",X"0D",X"20",X"09",X"FD",X"36",X"02",X"BB",
		X"DD",X"36",X"02",X"BC",X"C9",X"3A",X"26",X"F0",X"FE",X"01",X"C0",X"78",X"FE",X"07",X"20",X"09",
		X"FD",X"36",X"02",X"BD",X"DD",X"36",X"02",X"BE",X"C9",X"FE",X"01",X"C0",X"FD",X"36",X"00",X"00",
		X"DD",X"36",X"00",X"00",X"3A",X"AD",X"F0",X"D6",X"02",X"32",X"AD",X"F0",X"C9",X"E1",X"34",X"3E",
		X"02",X"32",X"09",X"F4",X"3A",X"7A",X"F3",X"B7",X"C2",X"43",X"6E",X"3A",X"89",X"F3",X"B7",X"20",
		X"31",X"32",X"12",X"F0",X"3A",X"60",X"F0",X"B7",X"28",X"12",X"AF",X"32",X"58",X"F0",X"DD",X"2A",
		X"5F",X"F0",X"DD",X"36",X"02",X"15",X"32",X"60",X"F0",X"32",X"58",X"F0",X"32",X"57",X"F0",X"32",
		X"5E",X"F0",X"32",X"43",X"F0",X"32",X"8A",X"F3",X"0E",X"01",X"CD",X"4E",X"3D",X"3E",X"80",X"C3",
		X"67",X"71",X"3D",X"32",X"89",X"F3",X"FE",X"08",X"30",X"09",X"ED",X"44",X"21",X"70",X"E8",X"85",
		X"6F",X"36",X"00",X"3A",X"0A",X"F0",X"B7",X"28",X"09",X"32",X"0C",X"F0",X"21",X"B0",X"F0",X"36",
		X"09",X"C9",X"3A",X"AE",X"F0",X"B7",X"28",X"0B",X"21",X"82",X"F0",X"36",X"04",X"21",X"B0",X"F0",
		X"36",X"0B",X"C9",X"3A",X"A0",X"F0",X"FE",X"01",X"20",X"12",X"AF",X"32",X"33",X"F0",X"32",X"35",
		X"F0",X"21",X"82",X"F0",X"36",X"04",X"21",X"B0",X"F0",X"36",X"0A",X"C9",X"FE",X"03",X"20",X"06",
		X"21",X"07",X"F0",X"4E",X"18",X"40",X"06",X"00",X"0E",X"F8",X"FD",X"21",X"5B",X"F2",X"CD",X"B5",
		X"41",X"3A",X"15",X"F0",X"B7",X"20",X"06",X"3A",X"AF",X"F0",X"B7",X"28",X"0B",X"FD",X"7E",X"02",
		X"B7",X"28",X"05",X"FD",X"7E",X"03",X"18",X"0A",X"FD",X"7E",X"01",X"FE",X"60",X"30",X"03",X"FD",
		X"7E",X"03",X"4F",X"3A",X"15",X"F0",X"B7",X"3E",X"D0",X"28",X"02",X"3E",X"E8",X"81",X"4F",X"3A",
		X"07",X"F0",X"B9",X"20",X"01",X"0D",X"DD",X"21",X"8B",X"F2",X"06",X"06",X"11",X"23",X"00",X"DD",
		X"7E",X"01",X"B7",X"28",X"1B",X"DD",X"19",X"10",X"F6",X"DD",X"21",X"8B",X"F2",X"06",X"06",X"DD",
		X"7E",X"05",X"B7",X"28",X"08",X"DD",X"19",X"10",X"F6",X"DD",X"21",X"8B",X"F2",X"CD",X"32",X"3F",
		X"21",X"32",X"F0",X"34",X"DD",X"22",X"B2",X"F0",X"DD",X"36",X"01",X"01",X"DD",X"71",X"05",X"DD",
		X"36",X"07",X"F8",X"3A",X"07",X"F0",X"B9",X"3E",X"00",X"20",X"01",X"3D",X"DD",X"77",X"08",X"DD",
		X"36",X"1E",X"00",X"3A",X"15",X"F0",X"B7",X"3E",X"29",X"28",X"02",X"3E",X"8A",X"DD",X"77",X"06",
		X"3C",X"DD",X"77",X"1D",X"3A",X"E6",X"BA",X"DD",X"77",X"0E",X"3A",X"EF",X"BA",X"DD",X"77",X"0F",
		X"DD",X"36",X"1F",X"00",X"DD",X"36",X"0A",X"00",X"3A",X"15",X"F0",X"B7",X"20",X"21",X"DD",X"36",
		X"02",X"15",X"DD",X"36",X"1C",X"06",X"DD",X"36",X"10",X"FD",X"3A",X"07",X"F0",X"DD",X"96",X"05",
		X"28",X"06",X"3E",X"01",X"30",X"02",X"ED",X"44",X"32",X"B1",X"F0",X"DD",X"77",X"04",X"C9",X"DD",
		X"36",X"02",X"95",X"DD",X"36",X"04",X"00",X"DD",X"36",X"10",X"FE",X"DD",X"36",X"01",X"01",X"3E",
		X"02",X"32",X"B1",X"F0",X"3A",X"03",X"F0",X"F6",X"20",X"32",X"03",X"F0",X"DD",X"21",X"6C",X"F8",
		X"DD",X"36",X"02",X"84",X"DD",X"36",X"06",X"85",X"0E",X"4F",X"CD",X"4E",X"3D",X"C9",X"DD",X"2A",
		X"B2",X"F0",X"3A",X"15",X"F0",X"B7",X"20",X"64",X"DD",X"7E",X"08",X"B7",X"28",X"13",X"DD",X"7E",
		X"07",X"C6",X"03",X"DD",X"77",X"07",X"E1",X"D0",X"AF",X"DD",X"77",X"08",X"32",X"07",X"F0",X"18",
		X"30",X"DD",X"7E",X"07",X"D6",X"03",X"DD",X"77",X"07",X"DD",X"35",X"1C",X"20",X"11",X"DD",X"36",
		X"1C",X"06",X"DD",X"7E",X"06",X"06",X"29",X"B8",X"20",X"02",X"06",X"D3",X"DD",X"70",X"06",X"3A",
		X"B1",X"F0",X"DD",X"77",X"04",X"DD",X"86",X"05",X"DD",X"77",X"05",X"21",X"07",X"F0",X"BE",X"E1",
		X"C0",X"34",X"DD",X"36",X"04",X"00",X"DD",X"7E",X"07",X"FE",X"A0",X"3E",X"00",X"28",X"06",X"3C",
		X"3C",X"38",X"02",X"ED",X"44",X"32",X"B1",X"F0",X"DD",X"77",X"10",X"C9",X"E1",X"23",X"DD",X"7E",
		X"07",X"96",X"DD",X"77",X"07",X"4F",X"06",X"00",X"FD",X"21",X"5B",X"F2",X"CD",X"B5",X"41",X"FD",
		X"7E",X"02",X"B7",X"28",X"05",X"FD",X"7E",X"03",X"18",X"0A",X"FD",X"7E",X"01",X"FE",X"60",X"30",
		X"03",X"FD",X"7E",X"03",X"C6",X"E8",X"DD",X"BE",X"05",X"28",X"0A",X"38",X"05",X"DD",X"34",X"05",
		X"18",X"03",X"DD",X"35",X"05",X"79",X"FE",X"D9",X"D0",X"FD",X"21",X"6C",X"F8",X"DD",X"46",X"05",
		X"FE",X"C9",X"30",X"09",X"FD",X"70",X"04",X"C6",X"30",X"FD",X"77",X"07",X"79",X"FD",X"70",X"00",
		X"C6",X"20",X"FD",X"77",X"03",X"32",X"01",X"F0",X"78",X"32",X"00",X"F0",X"32",X"07",X"F0",X"79",
		X"FE",X"C0",X"D0",X"FE",X"B0",X"28",X"0B",X"3E",X"01",X"32",X"B1",X"F0",X"ED",X"44",X"DD",X"77",
		X"10",X"C9",X"21",X"B0",X"F0",X"36",X"07",X"DD",X"36",X"03",X"02",X"DD",X"36",X"0B",X"04",X"DD",
		X"36",X"04",X"FF",X"C9",X"E1",X"FD",X"2A",X"B2",X"F0",X"FD",X"36",X"04",X"00",X"FD",X"35",X"1C",
		X"20",X"11",X"FD",X"36",X"1C",X"06",X"FD",X"7E",X"06",X"06",X"29",X"B8",X"20",X"02",X"06",X"D3",
		X"FD",X"70",X"06",X"3A",X"B1",X"F0",X"47",X"FD",X"86",X"07",X"FD",X"77",X"07",X"CB",X"78",X"28",
		X"05",X"FE",X"A2",X"38",X"04",X"C9",X"FE",X"A0",X"D8",X"FD",X"36",X"07",X"A0",X"FD",X"36",X"06",
		X"29",X"34",X"23",X"36",X"10",X"21",X"00",X"F0",X"FD",X"7E",X"05",X"77",X"23",X"36",X"AC",X"23",
		X"36",X"08",X"FD",X"21",X"68",X"F8",X"FD",X"77",X"00",X"FD",X"36",X"02",X"2B",X"FD",X"36",X"03",
		X"B0",X"C9",X"E1",X"FD",X"21",X"68",X"F8",X"FD",X"34",X"03",X"23",X"35",X"C0",X"2B",X"34",X"C9",
		X"E1",X"3A",X"01",X"F0",X"C6",X"02",X"32",X"01",X"F0",X"FE",X"D0",X"C0",X"34",X"21",X"68",X"F8",
		X"36",X"00",X"FD",X"2A",X"B2",X"F0",X"FD",X"36",X"03",X"04",X"FD",X"36",X"0B",X"06",X"FD",X"36",
		X"04",X"FE",X"3A",X"60",X"F0",X"B7",X"CC",X"6B",X"24",X"C9",X"DD",X"2A",X"B2",X"F0",X"DD",X"7E",
		X"07",X"D6",X"04",X"DD",X"77",X"07",X"CD",X"F3",X"43",X"DD",X"7E",X"05",X"DD",X"86",X"04",X"DD",
		X"77",X"05",X"47",X"FD",X"21",X"5B",X"F2",X"CD",X"62",X"45",X"E1",X"38",X"05",X"DD",X"36",X"04",
		X"FE",X"C9",X"DD",X"71",X"09",X"34",X"21",X"AF",X"F0",X"71",X"C9",X"DD",X"2A",X"B2",X"F0",X"DD",
		X"36",X"01",X"80",X"DD",X"36",X"0C",X"01",X"3A",X"01",X"F4",X"B7",X"3A",X"12",X"F0",X"20",X"02",
		X"F6",X"01",X"32",X"12",X"F0",X"AF",X"E1",X"36",X"00",X"32",X"03",X"F0",X"21",X"09",X"F4",X"36",
		X"01",X"3A",X"83",X"F0",X"EE",X"10",X"32",X"83",X"F0",X"21",X"05",X"F0",X"36",X"04",X"21",X"06",
		X"F0",X"36",X"02",X"3A",X"07",X"F0",X"B7",X"20",X"13",X"3A",X"00",X"F0",X"32",X"07",X"F0",X"3A",
		X"E5",X"F0",X"B7",X"C0",X"3C",X"32",X"E5",X"F0",X"32",X"E6",X"F0",X"C9",X"3A",X"36",X"F0",X"32",
		X"35",X"F0",X"3A",X"15",X"F0",X"B7",X"C8",X"21",X"38",X"F0",X"36",X"C0",X"C9",X"06",X"00",X"CD",
		X"CB",X"2B",X"CD",X"40",X"2C",X"3A",X"0A",X"F0",X"06",X"FF",X"FE",X"01",X"28",X"01",X"04",X"21",
		X"0D",X"F0",X"86",X"77",X"B8",X"E1",X"C0",X"36",X"03",X"AF",X"32",X"0A",X"F0",X"32",X"0C",X"F0",
		X"32",X"AF",X"F0",X"32",X"06",X"F0",X"C3",X"86",X"6E",X"06",X"00",X"0E",X"F0",X"FD",X"21",X"5B",
		X"F2",X"CD",X"B5",X"41",X"21",X"A0",X"F0",X"7E",X"FE",X"01",X"FD",X"7E",X"00",X"20",X"06",X"B7",
		X"20",X"01",X"34",X"E1",X"C9",X"B7",X"28",X"FB",X"34",X"E1",X"36",X"03",X"FD",X"7E",X"01",X"C6",
		X"03",X"32",X"07",X"F0",X"4F",X"AF",X"32",X"AF",X"F0",X"32",X"06",X"F0",X"32",X"82",X"F0",X"C3",
		X"C6",X"6E",X"E1",X"3A",X"AE",X"F0",X"B7",X"C0",X"36",X"03",X"AF",X"32",X"82",X"F0",X"C3",X"86",
		X"6E",X"3A",X"88",X"F0",X"B7",X"3E",X"20",X"28",X"02",X"3E",X"10",X"21",X"87",X"F0",X"96",X"80",
		X"CB",X"3F",X"E6",X"F0",X"47",X"3E",X"F0",X"91",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"B0",X"57",X"2A",X"91",X"F0",X"01",X"22",X"00",X"09",X"CB",X"2C",X"CB",X"1D",X"06",X"E0",X"0E",
		X"E3",X"3A",X"15",X"F0",X"B7",X"28",X"04",X"06",X"E4",X"0E",X"E7",X"7C",X"E6",X"03",X"80",X"67",
		X"7D",X"E6",X"F0",X"82",X"30",X"08",X"24",X"F5",X"7C",X"F6",X"E4",X"A1",X"67",X"F1",X"6F",X"C9",
		X"21",X"25",X"F0",X"36",X"01",X"DD",X"E5",X"DD",X"21",X"78",X"F8",X"DD",X"36",X"00",X"00",X"DD",
		X"36",X"04",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"0C",X"00",X"DD",X"36",X"10",X"00",X"DD",
		X"36",X"14",X"00",X"DD",X"E1",X"C9",X"3A",X"B8",X"F0",X"B7",X"28",X"08",X"3A",X"B9",X"F0",X"FE",
		X"06",X"DA",X"2D",X"73",X"3A",X"03",X"F0",X"E6",X"20",X"20",X"7F",X"16",X"00",X"3A",X"09",X"F0",
		X"B7",X"20",X"07",X"3A",X"06",X"F0",X"FE",X"02",X"20",X"0F",X"3A",X"82",X"F0",X"B7",X"28",X"09",
		X"3A",X"13",X"F0",X"57",X"ED",X"44",X"32",X"13",X"F0",X"21",X"67",X"B9",X"3A",X"15",X"F0",X"B7",
		X"28",X"03",X"21",X"9D",X"B9",X"3A",X"02",X"F0",X"CB",X"27",X"47",X"CB",X"27",X"80",X"85",X"30",
		X"01",X"24",X"6F",X"E5",X"FD",X"E1",X"DD",X"21",X"6C",X"F8",X"FD",X"7E",X"00",X"DD",X"77",X"02",
		X"3C",X"DD",X"77",X"06",X"FD",X"7E",X"01",X"DD",X"77",X"01",X"DD",X"77",X"05",X"3A",X"00",X"F0",
		X"FD",X"86",X"02",X"82",X"DD",X"77",X"00",X"3A",X"01",X"F0",X"FD",X"86",X"03",X"DD",X"77",X"03",
		X"3A",X"00",X"F0",X"FD",X"86",X"04",X"82",X"DD",X"77",X"04",X"3A",X"01",X"F0",X"FD",X"86",X"05",
		X"DD",X"77",X"07",X"CD",X"1C",X"75",X"3A",X"15",X"F0",X"B7",X"C4",X"41",X"75",X"DD",X"21",X"A8",
		X"F8",X"FD",X"21",X"8B",X"F2",X"01",X"04",X"00",X"2E",X"06",X"FD",X"7E",X"05",X"B7",X"CA",X"10",
		X"74",X"67",X"FD",X"7E",X"02",X"E6",X"10",X"20",X"59",X"DD",X"74",X"00",X"CD",X"7F",X"74",X"FD",
		X"7E",X"07",X"DD",X"77",X"03",X"DD",X"09",X"FD",X"7E",X"18",X"B7",X"20",X"06",X"CD",X"78",X"79",
		X"C3",X"73",X"74",X"57",X"FD",X"5E",X"17",X"FD",X"7E",X"19",X"FE",X"80",X"20",X"04",X"1A",X"3C",
		X"18",X"03",X"FD",X"86",X"05",X"12",X"13",X"AF",X"12",X"13",X"FD",X"7E",X"1B",X"12",X"13",X"FD",
		X"7E",X"07",X"FD",X"86",X"1A",X"67",X"FD",X"7E",X"08",X"B7",X"7C",X"28",X"06",X"FE",X"F7",X"30",
		X"0D",X"18",X"04",X"FE",X"F7",X"38",X"07",X"AF",X"12",X"1B",X"12",X"1B",X"12",X"1B",X"12",X"C3",
		X"73",X"74",X"3A",X"15",X"F0",X"B7",X"28",X"06",X"CD",X"71",X"78",X"CD",X"E6",X"77",X"FD",X"7E",
		X"08",X"B7",X"20",X"27",X"DD",X"74",X"00",X"FD",X"56",X"06",X"DD",X"72",X"02",X"FD",X"7E",X"07",
		X"DD",X"77",X"03",X"DD",X"09",X"FE",X"E7",X"30",X"65",X"C6",X"10",X"DD",X"77",X"03",X"7C",X"FD",
		X"86",X"1E",X"DD",X"77",X"00",X"CD",X"BB",X"74",X"C3",X"57",X"73",X"FD",X"7E",X"07",X"FE",X"F7",
		X"30",X"0E",X"DD",X"36",X"00",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"00",X"18",X"0C",
		X"DD",X"74",X"00",X"FD",X"56",X"06",X"DD",X"72",X"02",X"DD",X"77",X"03",X"DD",X"09",X"C6",X"10",
		X"DD",X"77",X"03",X"7C",X"FD",X"86",X"1E",X"DD",X"77",X"00",X"CD",X"BB",X"74",X"C3",X"57",X"73",
		X"DD",X"77",X"00",X"DD",X"77",X"02",X"DD",X"77",X"03",X"FD",X"7E",X"09",X"FE",X"03",X"20",X"0C",
		X"11",X"F4",X"F8",X"AF",X"12",X"11",X"F8",X"F8",X"12",X"FD",X"77",X"09",X"DD",X"09",X"DD",X"36",
		X"00",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"00",X"FD",X"7E",X"09",X"FE",X"03",X"20",
		X"05",X"11",X"F8",X"F8",X"AF",X"12",X"FD",X"7E",X"18",X"B7",X"28",X"09",X"57",X"FD",X"5E",X"17",
		X"AF",X"12",X"FD",X"77",X"18",X"FD",X"7E",X"13",X"B7",X"28",X"09",X"57",X"FD",X"5E",X"12",X"AF",
		X"12",X"FD",X"77",X"13",X"FD",X"7E",X"15",X"B7",X"28",X"09",X"57",X"FD",X"5E",X"14",X"AF",X"12",
		X"FD",X"77",X"15",X"DD",X"09",X"11",X"23",X"00",X"FD",X"19",X"2D",X"C2",X"3A",X"73",X"C9",X"FD",
		X"56",X"06",X"FD",X"7E",X"01",X"E6",X"0F",X"20",X"2E",X"FD",X"7E",X"08",X"B7",X"20",X"28",X"FD",
		X"7E",X"10",X"CB",X"7F",X"20",X"21",X"B7",X"28",X"1E",X"FD",X"35",X"22",X"C0",X"FD",X"36",X"22",
		X"01",X"FD",X"7E",X"21",X"EE",X"01",X"FD",X"77",X"21",X"28",X"0C",X"FD",X"7E",X"02",X"E6",X"0F",
		X"FE",X"02",X"16",X"78",X"28",X"01",X"15",X"DD",X"72",X"02",X"C9",X"FD",X"56",X"1D",X"3A",X"15",
		X"F0",X"B7",X"20",X"54",X"FD",X"7E",X"01",X"E6",X"0F",X"20",X"4D",X"FD",X"7E",X"08",X"B7",X"20",
		X"47",X"FD",X"7E",X"10",X"CB",X"7F",X"20",X"40",X"B7",X"28",X"3D",X"FD",X"7E",X"02",X"E6",X"0F",
		X"FE",X"04",X"28",X"09",X"30",X"32",X"FD",X"7E",X"10",X"FE",X"06",X"38",X"2B",X"FD",X"35",X"22",
		X"C0",X"FD",X"36",X"22",X"01",X"FD",X"7E",X"21",X"EE",X"01",X"FD",X"77",X"21",X"28",X"19",X"FD",
		X"7E",X"02",X"E6",X"0F",X"16",X"79",X"28",X"10",X"FE",X"04",X"16",X"88",X"28",X"0A",X"14",X"FD",
		X"7E",X"1D",X"FE",X"7D",X"28",X"02",X"16",X"7A",X"DD",X"72",X"02",X"C9",X"3A",X"D5",X"F0",X"B7",
		X"C0",X"3A",X"24",X"F0",X"B7",X"C8",X"FE",X"03",X"D0",X"C6",X"12",X"21",X"01",X"F0",X"86",X"DD",
		X"21",X"FC",X"F8",X"DD",X"77",X"03",X"3A",X"00",X"F0",X"FD",X"86",X"04",X"82",X"DD",X"77",X"00",
		X"C9",X"3A",X"03",X"F0",X"47",X"E6",X"40",X"28",X"06",X"CD",X"92",X"76",X"C3",X"6A",X"76",X"0E",
		X"04",X"3A",X"FF",X"F0",X"B7",X"28",X"06",X"FE",X"03",X"30",X"02",X"0E",X"F4",X"78",X"E6",X"20",
		X"20",X"12",X"0D",X"3A",X"82",X"F0",X"FE",X"0A",X"30",X"0A",X"0D",X"FE",X"06",X"30",X"05",X"0D",
		X"B7",X"20",X"01",X"0D",X"3A",X"20",X"F0",X"B9",X"28",X"0E",X"AF",X"32",X"1B",X"F0",X"3C",X"32",
		X"1D",X"F0",X"79",X"32",X"20",X"F0",X"18",X"05",X"E6",X"0F",X"CA",X"6A",X"76",X"DD",X"21",X"48",
		X"F8",X"21",X"1D",X"F0",X"35",X"20",X"36",X"36",X"04",X"3A",X"1B",X"F0",X"3C",X"FE",X"06",X"38",
		X"01",X"AF",X"32",X"1B",X"F0",X"21",X"F3",X"BB",X"CB",X"27",X"85",X"30",X"01",X"24",X"6F",X"5E",
		X"23",X"56",X"D5",X"E1",X"11",X"04",X"00",X"06",X"06",X"CB",X"79",X"28",X"02",X"06",X"04",X"7E",
		X"DD",X"77",X"02",X"23",X"7E",X"DD",X"77",X"01",X"23",X"DD",X"19",X"10",X"F2",X"79",X"E6",X"0F",
		X"6F",X"CB",X"27",X"85",X"21",X"F2",X"75",X"85",X"30",X"01",X"24",X"6F",X"DD",X"21",X"48",X"F8",
		X"11",X"04",X"00",X"3A",X"00",X"F0",X"C6",X"08",X"47",X"D6",X"10",X"4F",X"3A",X"01",X"F0",X"C6",
		X"06",X"E9",X"C3",X"01",X"76",X"C3",X"1A",X"76",X"C3",X"2E",X"76",X"C3",X"49",X"76",X"C3",X"1A",
		X"76",X"06",X"06",X"3A",X"20",X"F0",X"CB",X"7F",X"28",X"05",X"05",X"05",X"CA",X"6A",X"76",X"DD",
		X"36",X"00",X"00",X"DD",X"19",X"10",X"F8",X"C3",X"6A",X"76",X"DD",X"70",X"00",X"DD",X"77",X"03",
		X"DD",X"19",X"DD",X"71",X"00",X"DD",X"77",X"03",X"DD",X"19",X"06",X"04",X"18",X"D5",X"26",X"02",
		X"DD",X"70",X"00",X"DD",X"77",X"03",X"DD",X"19",X"DD",X"71",X"00",X"DD",X"77",X"03",X"DD",X"19",
		X"C6",X"10",X"25",X"20",X"EB",X"06",X"02",X"18",X"BA",X"F5",X"26",X"03",X"3A",X"20",X"F0",X"CB",
		X"7F",X"28",X"01",X"25",X"F1",X"DD",X"70",X"00",X"DD",X"77",X"03",X"DD",X"19",X"DD",X"71",X"00",
		X"DD",X"77",X"03",X"DD",X"19",X"C6",X"10",X"25",X"20",X"EB",X"3A",X"7E",X"F0",X"B7",X"C8",X"06",
		X"00",X"FE",X"10",X"38",X"01",X"04",X"3A",X"21",X"F0",X"3C",X"32",X"21",X"F0",X"CB",X"57",X"28",
		X"02",X"06",X"02",X"DD",X"21",X"70",X"F8",X"DD",X"7E",X"02",X"FE",X"85",X"C0",X"80",X"DD",X"77",
		X"02",X"C9",X"3A",X"22",X"F0",X"47",X"CB",X"27",X"80",X"21",X"A9",X"76",X"85",X"30",X"01",X"24",
		X"6F",X"11",X"04",X"00",X"DD",X"21",X"48",X"F8",X"E9",X"C3",X"C1",X"76",X"C3",X"14",X"77",X"C3",
		X"37",X"77",X"C3",X"91",X"77",X"C3",X"91",X"77",X"C3",X"91",X"77",X"C3",X"91",X"77",X"C3",X"C6",
		X"77",X"3A",X"82",X"F0",X"CB",X"3F",X"FE",X"08",X"38",X"02",X"3E",X"07",X"32",X"23",X"F0",X"47",
		X"21",X"00",X"F0",X"86",X"DD",X"77",X"00",X"3A",X"01",X"F0",X"C6",X"0A",X"CB",X"38",X"80",X"DD",
		X"77",X"03",X"DD",X"36",X"02",X"31",X"DD",X"36",X"01",X"00",X"06",X"05",X"3A",X"FF",X"F0",X"B7",
		X"28",X"06",X"FE",X"03",X"30",X"02",X"06",X"03",X"DD",X"19",X"DD",X"36",X"00",X"00",X"10",X"F8",
		X"DD",X"21",X"6C",X"F8",X"DD",X"36",X"02",X"D4",X"DD",X"36",X"06",X"D5",X"3E",X"09",X"32",X"02",
		X"F0",X"C3",X"E1",X"77",X"3A",X"23",X"F0",X"B7",X"28",X"18",X"3D",X"32",X"23",X"F0",X"47",X"21",
		X"00",X"F0",X"86",X"DD",X"77",X"00",X"3A",X"01",X"F0",X"C6",X"0A",X"CB",X"38",X"80",X"DD",X"77",
		X"03",X"C9",X"3E",X"08",X"32",X"02",X"F0",X"0E",X"33",X"CD",X"4E",X"3D",X"3A",X"00",X"F0",X"C6",
		X"08",X"DD",X"77",X"00",X"47",X"3A",X"01",X"F0",X"D6",X"04",X"DD",X"77",X"03",X"4F",X"DD",X"36",
		X"02",X"64",X"DD",X"36",X"01",X"00",X"DD",X"19",X"78",X"D6",X"10",X"67",X"DD",X"77",X"00",X"DD",
		X"71",X"03",X"DD",X"36",X"02",X"66",X"DD",X"36",X"01",X"00",X"DD",X"19",X"DD",X"74",X"00",X"79",
		X"C6",X"10",X"4F",X"DD",X"77",X"03",X"DD",X"36",X"02",X"67",X"DD",X"36",X"01",X"00",X"DD",X"19",
		X"DD",X"70",X"00",X"DD",X"71",X"03",X"DD",X"36",X"02",X"65",X"DD",X"36",X"01",X"00",X"C3",X"E1",
		X"77",X"3A",X"00",X"F0",X"C6",X"08",X"DD",X"77",X"00",X"47",X"3A",X"01",X"F0",X"D6",X"04",X"DD",
		X"77",X"03",X"4F",X"DD",X"19",X"78",X"D6",X"10",X"67",X"DD",X"77",X"00",X"DD",X"71",X"03",X"DD",
		X"19",X"DD",X"74",X"00",X"79",X"C6",X"10",X"4F",X"DD",X"77",X"03",X"DD",X"19",X"DD",X"70",X"00",
		X"DD",X"71",X"03",X"C3",X"E1",X"77",X"AF",X"06",X"04",X"DD",X"77",X"00",X"DD",X"19",X"10",X"F9",
		X"32",X"22",X"F0",X"3A",X"03",X"F0",X"EE",X"40",X"32",X"03",X"F0",X"21",X"20",X"F0",X"36",X"FF",
		X"C9",X"21",X"22",X"F0",X"34",X"C9",X"FD",X"7E",X"06",X"FE",X"8A",X"C0",X"FD",X"7E",X"08",X"B7",
		X"C0",X"FD",X"7E",X"07",X"FE",X"E7",X"D0",X"FD",X"7E",X"01",X"E6",X"0A",X"C0",X"FD",X"7E",X"18",
		X"B7",X"20",X"1F",X"FD",X"E5",X"CD",X"EF",X"1B",X"30",X"06",X"01",X"04",X"00",X"FD",X"E1",X"C9",
		X"FD",X"E5",X"C1",X"FD",X"E1",X"FD",X"71",X"17",X"FD",X"70",X"18",X"01",X"04",X"00",X"FD",X"36",
		X"1C",X"00",X"FD",X"7E",X"1C",X"B7",X"20",X"0E",X"FD",X"36",X"1B",X"8C",X"FD",X"36",X"19",X"00",
		X"FD",X"36",X"1A",X"0A",X"18",X"34",X"FE",X"04",X"38",X"30",X"20",X"06",X"FD",X"36",X"1B",X"8D",
		X"18",X"28",X"FE",X"08",X"38",X"24",X"20",X"0E",X"FD",X"36",X"1B",X"8E",X"FD",X"36",X"19",X"80",
		X"FD",X"36",X"1A",X"10",X"18",X"14",X"FE",X"0C",X"20",X"04",X"FD",X"36",X"1B",X"8F",X"FD",X"7E",
		X"1A",X"FD",X"86",X"03",X"FD",X"77",X"1A",X"FD",X"7E",X"1C",X"3C",X"E6",X"0F",X"FD",X"77",X"1C",
		X"C9",X"FD",X"7E",X"02",X"E6",X"80",X"C8",X"FD",X"7E",X"08",X"FE",X"01",X"38",X"1F",X"C8",X"FD",
		X"7E",X"07",X"FE",X"F7",X"30",X"1D",X"FD",X"7E",X"13",X"B7",X"C8",X"57",X"FD",X"5E",X"12",X"AF",
		X"12",X"FD",X"7E",X"15",X"B7",X"C8",X"57",X"FD",X"5E",X"14",X"AF",X"12",X"C9",X"FD",X"7E",X"07",
		X"FE",X"E7",X"D0",X"E5",X"DD",X"E5",X"FD",X"E5",X"DD",X"E1",X"6F",X"DD",X"66",X"05",X"DD",X"7E",
		X"13",X"B7",X"20",X"2B",X"CD",X"CD",X"40",X"30",X"0B",X"01",X"04",X"00",X"DD",X"E5",X"FD",X"E1",
		X"DD",X"E1",X"E1",X"C9",X"FD",X"36",X"02",X"AF",X"FD",X"36",X"01",X"00",X"FD",X"E5",X"C1",X"DD",
		X"71",X"12",X"DD",X"70",X"13",X"DD",X"36",X"21",X"00",X"DD",X"36",X"22",X"04",X"18",X"09",X"DD",
		X"4E",X"12",X"DD",X"46",X"13",X"C5",X"FD",X"E1",X"06",X"03",X"0E",X"0D",X"DD",X"7E",X"02",X"E6",
		X"0F",X"FE",X"01",X"28",X"04",X"06",X"04",X"0E",X"11",X"7C",X"80",X"FD",X"77",X"00",X"7C",X"90",
		X"67",X"7D",X"81",X"FD",X"77",X"03",X"6F",X"DD",X"35",X"22",X"20",X"15",X"DD",X"36",X"22",X"04",
		X"DD",X"7E",X"21",X"EE",X"01",X"DD",X"77",X"21",X"06",X"AF",X"28",X"02",X"06",X"B3",X"FD",X"70",
		X"02",X"DD",X"7E",X"15",X"B7",X"20",X"23",X"CD",X"CD",X"40",X"30",X"0B",X"01",X"04",X"00",X"DD",
		X"E5",X"FD",X"E1",X"DD",X"E1",X"E1",X"C9",X"FD",X"36",X"02",X"AF",X"FD",X"36",X"01",X"20",X"FD",
		X"E5",X"C1",X"DD",X"71",X"14",X"DD",X"70",X"15",X"18",X"09",X"DD",X"4E",X"14",X"DD",X"46",X"15",
		X"C5",X"FD",X"E1",X"FD",X"74",X"00",X"FD",X"75",X"03",X"DD",X"7E",X"22",X"FE",X"04",X"20",X"0D",
		X"DD",X"7E",X"21",X"B7",X"06",X"AF",X"28",X"02",X"06",X"B3",X"FD",X"70",X"02",X"DD",X"E5",X"FD",
		X"E1",X"DD",X"E1",X"E1",X"01",X"04",X"00",X"C9",X"FD",X"7E",X"02",X"E6",X"80",X"C8",X"FD",X"7E",
		X"01",X"E6",X"0A",X"C0",X"FD",X"E5",X"CD",X"EF",X"1B",X"01",X"04",X"00",X"30",X"03",X"FD",X"E1",
		X"C9",X"FD",X"E5",X"D1",X"FD",X"E1",X"FD",X"72",X"18",X"FD",X"73",X"17",X"FD",X"36",X"1A",X"07",
		X"FD",X"7E",X"02",X"E6",X"01",X"FD",X"77",X"19",X"3E",X"AD",X"28",X"02",X"3E",X"74",X"FD",X"77",
		X"1B",X"F1",X"C3",X"57",X"73",X"3A",X"03",X"F0",X"47",X"E6",X"10",X"C0",X"3A",X"15",X"F0",X"21",
		X"16",X"F0",X"BE",X"C0",X"3A",X"0A",X"F0",X"FE",X"01",X"38",X"79",X"C0",X"78",X"E6",X"41",X"C0",
		X"21",X"01",X"F0",X"1E",X"00",X"16",X"00",X"3E",X"D0",X"96",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"47",X"21",X"5D",X"7F",X"3A",X"0B",X"F0",X"80",X"D6",X"46",X"38",X"0D",X"FE",X"3B",
		X"38",X"02",X"3E",X"3B",X"5F",X"85",X"30",X"01",X"24",X"6F",X"14",X"3A",X"0D",X"F0",X"86",X"FE",
		X"60",X"30",X"02",X"3E",X"FF",X"4F",X"21",X"00",X"F0",X"96",X"30",X"21",X"7B",X"B7",X"20",X"2C",
		X"3A",X"A1",X"F0",X"CB",X"7F",X"C8",X"71",X"0E",X"12",X"CD",X"4E",X"3D",X"3E",X"04",X"32",X"A1",
		X"F0",X"32",X"27",X"F0",X"3A",X"03",X"F0",X"F6",X"04",X"32",X"03",X"F0",X"C9",X"FE",X"14",X"D0",
		X"7A",X"B7",X"C8",X"3A",X"03",X"F0",X"F6",X"40",X"32",X"03",X"F0",X"C9",X"3E",X"FE",X"32",X"A1",
		X"F0",X"C3",X"AF",X"7D",X"CD",X"8F",X"1D",X"D2",X"A2",X"7D",X"3A",X"06",X"F0",X"FE",X"02",X"CA",
		X"F7",X"7C",X"1E",X"00",X"FD",X"21",X"8B",X"F2",X"FD",X"7E",X"01",X"E6",X"80",X"28",X"3D",X"FD",
		X"7E",X"05",X"B7",X"28",X"37",X"21",X"00",X"F0",X"47",X"FD",X"7E",X"02",X"E6",X"0F",X"FE",X"02",
		X"0E",X"02",X"38",X"02",X"0E",X"04",X"78",X"C6",X"10",X"91",X"BE",X"38",X"1F",X"7E",X"C6",X"10",
		X"91",X"B8",X"38",X"18",X"21",X"01",X"F0",X"FD",X"7E",X"07",X"47",X"FD",X"86",X"0E",X"D6",X"04",
		X"BE",X"38",X"09",X"3A",X"04",X"F0",X"D6",X"04",X"86",X"B8",X"30",X"0E",X"01",X"23",X"00",X"FD",
		X"09",X"1C",X"7B",X"FE",X"06",X"20",X"B1",X"C3",X"F7",X"7C",X"FD",X"7E",X"02",X"E6",X"0F",X"FE",
		X"06",X"38",X"17",X"3A",X"58",X"F0",X"FE",X"02",X"38",X"10",X"3A",X"00",X"F0",X"FD",X"96",X"05",
		X"CB",X"7F",X"28",X"02",X"ED",X"44",X"FE",X"03",X"38",X"D2",X"B7",X"20",X"0C",X"3A",X"A1",X"F0",
		X"CB",X"2F",X"CB",X"2F",X"FD",X"77",X"04",X"18",X"41",X"FD",X"7E",X"01",X"E6",X"40",X"28",X"3A",
		X"3A",X"01",X"F0",X"FD",X"96",X"07",X"30",X"02",X"ED",X"44",X"FE",X"0A",X"30",X"2C",X"3A",X"00",
		X"F0",X"FD",X"BE",X"05",X"30",X"0D",X"FD",X"7E",X"13",X"B7",X"28",X"1E",X"0E",X"F0",X"21",X"42",
		X"65",X"18",X"0B",X"FD",X"7E",X"15",X"B7",X"28",X"11",X"0E",X"10",X"21",X"16",X"65",X"FD",X"7E",
		X"05",X"81",X"32",X"00",X"F0",X"FD",X"E5",X"DD",X"E1",X"E9",X"0E",X"12",X"CD",X"4E",X"3D",X"FD",
		X"56",X"0F",X"26",X"03",X"3A",X"82",X"F0",X"6F",X"FD",X"7E",X"03",X"CD",X"22",X"7F",X"FD",X"66",
		X"0F",X"16",X"03",X"FD",X"6E",X"03",X"F5",X"3A",X"82",X"F0",X"CD",X"22",X"7F",X"CB",X"7F",X"28",
		X"05",X"FD",X"7E",X"03",X"CB",X"3F",X"FE",X"10",X"38",X"02",X"3E",X"0F",X"FD",X"77",X"03",X"FD",
		X"36",X"0D",X"04",X"3A",X"01",X"F0",X"47",X"C6",X"12",X"FD",X"96",X"07",X"30",X"16",X"FD",X"7E",
		X"07",X"C6",X"08",X"FD",X"77",X"07",X"3A",X"A1",X"F0",X"FD",X"B6",X"04",X"20",X"22",X"FD",X"36",
		X"04",X"02",X"18",X"1C",X"FD",X"7E",X"07",X"FD",X"86",X"0E",X"D6",X"04",X"B8",X"38",X"11",X"3A",
		X"00",X"F0",X"47",X"FD",X"BE",X"05",X"3E",X"0F",X"38",X"02",X"ED",X"44",X"80",X"FD",X"77",X"05",
		X"F1",X"CB",X"7F",X"28",X"05",X"3A",X"82",X"F0",X"CB",X"3F",X"FE",X"10",X"38",X"02",X"3E",X"0F",
		X"67",X"3A",X"03",X"F0",X"E6",X"01",X"20",X"13",X"2E",X"00",X"22",X"81",X"F0",X"CB",X"24",X"3A",
		X"84",X"F0",X"FE",X"10",X"20",X"02",X"CB",X"24",X"22",X"7F",X"F0",X"FD",X"56",X"0F",X"26",X"03",
		X"3A",X"A1",X"F0",X"ED",X"44",X"6F",X"FD",X"7E",X"04",X"CD",X"22",X"7F",X"FD",X"66",X"0F",X"16",
		X"03",X"FD",X"6E",X"04",X"F5",X"3A",X"A1",X"F0",X"ED",X"44",X"CD",X"22",X"7F",X"CD",X"51",X"7F",
		X"FD",X"77",X"04",X"3A",X"14",X"F0",X"B7",X"3E",X"05",X"28",X"02",X"CB",X"27",X"FD",X"86",X"0C",
		X"FD",X"77",X"0C",X"3E",X"03",X"BC",X"30",X"11",X"3A",X"00",X"F0",X"FD",X"BE",X"05",X"3E",X"08",
		X"30",X"02",X"ED",X"44",X"21",X"00",X"F0",X"86",X"77",X"C1",X"3A",X"03",X"F0",X"E6",X"02",X"20",
		X"0D",X"FD",X"7E",X"10",X"CB",X"7F",X"28",X"02",X"ED",X"44",X"FE",X"07",X"38",X"57",X"FD",X"7E",
		X"02",X"E6",X"0F",X"FE",X"06",X"30",X"3C",X"FD",X"7E",X"01",X"47",X"E6",X"08",X"28",X"14",X"78",
		X"EE",X"08",X"47",X"FD",X"7E",X"18",X"B7",X"28",X"0A",X"67",X"FD",X"6E",X"17",X"36",X"00",X"FD",
		X"36",X"18",X"00",X"FD",X"7E",X"1F",X"B7",X"20",X"17",X"78",X"F6",X"03",X"47",X"FD",X"36",X"1F",
		X"10",X"3A",X"01",X"F0",X"FD",X"BE",X"07",X"3E",X"01",X"38",X"02",X"C6",X"03",X"FD",X"77",X"03",
		X"FD",X"70",X"01",X"3A",X"03",X"F0",X"F6",X"02",X"32",X"03",X"F0",X"AF",X"32",X"A1",X"F0",X"3A",
		X"06",X"F0",X"C3",X"E7",X"7D",X"78",X"ED",X"44",X"CD",X"51",X"7F",X"32",X"A1",X"F0",X"CB",X"7F",
		X"28",X"02",X"ED",X"44",X"3C",X"32",X"27",X"F0",X"3A",X"03",X"F0",X"F6",X"04",X"32",X"03",X"F0",
		X"FD",X"7E",X"02",X"E6",X"0F",X"FE",X"06",X"38",X"11",X"3A",X"00",X"F0",X"FD",X"BE",X"05",X"3E",
		X"20",X"38",X"02",X"ED",X"44",X"FD",X"77",X"11",X"18",X"4D",X"06",X"04",X"FE",X"02",X"20",X"40",
		X"FD",X"7E",X"01",X"E6",X"0A",X"20",X"40",X"06",X"0A",X"FD",X"36",X"16",X"00",X"FD",X"36",X"20",
		X"18",X"FD",X"7E",X"04",X"B7",X"20",X"04",X"FD",X"36",X"04",X"02",X"21",X"28",X"F0",X"3A",X"8E",
		X"F3",X"3C",X"CB",X"27",X"C6",X"08",X"86",X"77",X"3A",X"5E",X"F0",X"B7",X"28",X"12",X"AF",X"32",
		X"5E",X"F0",X"3A",X"5D",X"F0",X"B7",X"20",X"08",X"3A",X"12",X"F0",X"EE",X"04",X"32",X"12",X"F0",
		X"FD",X"7E",X"01",X"B0",X"FD",X"77",X"01",X"3A",X"15",X"F0",X"B7",X"C2",X"BF",X"7E",X"06",X"02",
		X"11",X"04",X"00",X"FD",X"21",X"60",X"F8",X"DD",X"21",X"53",X"F0",X"21",X"00",X"F0",X"FD",X"7E",
		X"00",X"B7",X"28",X"58",X"4F",X"DD",X"7E",X"00",X"FE",X"10",X"79",X"20",X"08",X"C6",X"10",X"38",
		X"0A",X"BE",X"30",X"07",X"C9",X"D6",X"10",X"38",X"02",X"BE",X"D0",X"FD",X"36",X"00",X"00",X"3A",
		X"06",X"F0",X"FE",X"02",X"20",X"0D",X"3A",X"2F",X"F0",X"FE",X"04",X"30",X"18",X"3C",X"32",X"2F",
		X"F0",X"18",X"23",X"3A",X"01",X"F4",X"B7",X"28",X"0C",X"3A",X"2F",X"F0",X"B7",X"20",X"06",X"3C",
		X"32",X"2F",X"F0",X"18",X"11",X"3A",X"01",X"F0",X"C6",X"03",X"FD",X"BE",X"03",X"30",X"07",X"C6",
		X"08",X"FD",X"BE",X"03",X"30",X"0B",X"0E",X"37",X"CD",X"4E",X"3D",X"C9",X"FD",X"19",X"10",X"9E",
		X"C9",X"3A",X"42",X"F0",X"B7",X"28",X"07",X"3A",X"82",X"F0",X"FE",X"09",X"30",X"E8",X"3A",X"03",
		X"F0",X"F6",X"0A",X"32",X"03",X"F0",X"DD",X"7E",X"00",X"FE",X"10",X"3E",X"02",X"06",X"07",X"28",
		X"04",X"ED",X"44",X"06",X"00",X"32",X"A1",X"F0",X"21",X"02",X"F0",X"70",X"0E",X"35",X"CD",X"4E",
		X"3D",X"C9",X"3A",X"03",X"F0",X"47",X"E6",X"01",X"C2",X"52",X"7A",X"78",X"E6",X"40",X"C0",X"3A",
		X"06",X"F0",X"FE",X"02",X"38",X"31",X"3A",X"03",X"F0",X"E6",X"08",X"20",X"2D",X"3A",X"07",X"F0",
		X"21",X"00",X"F0",X"BE",X"30",X"01",X"77",X"CD",X"F7",X"7C",X"C9",X"3A",X"06",X"F0",X"FE",X"02",
		X"38",X"15",X"3A",X"00",X"F0",X"D6",X"20",X"32",X"00",X"F0",X"CD",X"8F",X"1D",X"3A",X"00",X"F0",
		X"C6",X"20",X"32",X"00",X"F0",X"18",X"E4",X"32",X"AF",X"F0",X"3A",X"19",X"F0",X"21",X"18",X"F0",
		X"B6",X"C0",X"3A",X"03",X"F0",X"47",X"E6",X"02",X"20",X"1A",X"3A",X"56",X"F0",X"FE",X"8E",X"28",
		X"13",X"21",X"A1",X"F0",X"7E",X"B7",X"20",X"03",X"3A",X"00",X"F0",X"FE",X"80",X"3E",X"02",X"30",
		X"02",X"ED",X"44",X"77",X"78",X"F6",X"03",X"32",X"03",X"F0",X"3A",X"B0",X"F0",X"B7",X"C0",X"CD",
		X"B3",X"3D",X"CD",X"E4",X"3D",X"3A",X"00",X"F0",X"FD",X"77",X"00",X"FD",X"36",X"01",X"00",X"3A",
		X"15",X"F0",X"B7",X"3E",X"21",X"28",X"02",X"3E",X"84",X"FD",X"77",X"02",X"3A",X"01",X"F0",X"FD",
		X"77",X"03",X"36",X"06",X"FD",X"22",X"2A",X"F0",X"CD",X"B3",X"3D",X"CD",X"E4",X"3D",X"3A",X"00",
		X"F0",X"FD",X"77",X"00",X"FD",X"36",X"01",X"00",X"3A",X"15",X"F0",X"B7",X"3E",X"22",X"28",X"02",
		X"3E",X"85",X"FD",X"77",X"02",X"3A",X"01",X"F0",X"C6",X"10",X"FD",X"77",X"03",X"36",X"06",X"FD",
		X"22",X"2C",X"F0",X"21",X"A6",X"F0",X"36",X"10",X"3A",X"35",X"F0",X"32",X"36",X"F0",X"AF",X"32",
		X"35",X"F0",X"32",X"45",X"F0",X"32",X"00",X"F0",X"32",X"01",X"F0",X"32",X"81",X"F0",X"32",X"82",
		X"F0",X"32",X"7F",X"F0",X"32",X"80",X"F0",X"32",X"D4",X"F0",X"32",X"FE",X"F0",X"3A",X"12",X"F0",
		X"E6",X"04",X"32",X"12",X"F0",X"CD",X"A0",X"52",X"3A",X"15",X"F0",X"B7",X"28",X"06",X"0E",X"12",
		X"CD",X"4E",X"3D",X"C9",X"3A",X"60",X"F0",X"B7",X"C8",X"21",X"5B",X"F0",X"36",X"02",X"C9",X"3A",
		X"C2",X"F0",X"B7",X"C8",X"FD",X"21",X"60",X"F8",X"06",X"02",X"21",X"C8",X"F0",X"FD",X"7E",X"00",
		X"B7",X"28",X"44",X"C6",X"08",X"4F",X"7E",X"FE",X"FF",X"28",X"3C",X"3A",X"00",X"F0",X"C6",X"08",
		X"91",X"30",X"02",X"ED",X"44",X"FE",X"07",X"30",X"2E",X"FD",X"7E",X"03",X"86",X"4F",X"3A",X"01",
		X"F0",X"C6",X"0C",X"91",X"30",X"02",X"ED",X"44",X"FE",X"0B",X"30",X"1B",X"FD",X"36",X"02",X"39",
		X"36",X"FF",X"23",X"36",X"06",X"0E",X"4C",X"3A",X"C2",X"F0",X"FE",X"02",X"DC",X"4E",X"3D",X"0E",
		X"13",X"CD",X"4E",X"3D",X"C3",X"AF",X"7D",X"05",X"C8",X"FD",X"21",X"64",X"F8",X"21",X"CA",X"F0",
		X"18",X"AB",X"CB",X"27",X"95",X"4F",X"42",X"AF",X"81",X"10",X"FD",X"5F",X"4D",X"44",X"AF",X"81",
		X"10",X"FD",X"83",X"5F",X"7C",X"82",X"47",X"7B",X"1E",X"00",X"CB",X"7F",X"28",X"04",X"1E",X"01",
		X"ED",X"44",X"0E",X"00",X"90",X"38",X"03",X"0C",X"18",X"FA",X"79",X"CB",X"43",X"C8",X"ED",X"44",
		X"C9",X"CB",X"7F",X"28",X"02",X"3C",X"C9",X"3D",X"CB",X"7F",X"C8",X"AF",X"C9",X"6D",X"50",X"3F",
		X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"3B",X"31",X"2B",X"2B",X"2B",X"2B",X"2B",X"26",X"1C",X"1C",
		X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"1C",X"0A",X"0A",X"0A",X"0A",X"0A",X"06",X"04",X"F9",X"F8",
		X"F8",X"F8",X"F8",X"F8",X"EC",X"EC",X"EC",X"E1",X"DA",X"DA",X"DA",X"D2",X"C9",X"BF",X"B9",X"B8",
		X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B8",X"B3",X"A9",X"16",X"00",X"DD",X"21",X"8B",X"F2",X"DD",
		X"7E",X"01",X"E6",X"80",X"CA",X"6C",X"83",X"DD",X"7E",X"05",X"B7",X"CA",X"6C",X"83",X"DD",X"7E",
		X"08",X"B7",X"C2",X"6C",X"83",X"DD",X"7E",X"1F",X"FE",X"0F",X"D2",X"6C",X"83",X"47",X"CB",X"27",
		X"80",X"21",X"CA",X"7F",X"85",X"30",X"01",X"24",X"6F",X"E9",X"C3",X"F7",X"7F",X"C3",X"38",X"81",
		X"C3",X"38",X"81",X"C3",X"38",X"81",X"C3",X"38",X"81",X"C3",X"3E",X"81",X"C3",X"CE",X"81",X"C3",
		X"CE",X"81",X"C3",X"CE",X"81",X"C3",X"32",X"3F",X"C3",X"38",X"81",X"C3",X"38",X"81",X"C3",X"38",
		X"81",X"C3",X"38",X"81",X"C3",X"B8",X"81",X"CD",X"30",X"20",X"DA",X"FA",X"81",X"DD",X"7E",X"01",
		X"47",X"E6",X"01",X"C2",X"FA",X"81",X"78",X"F6",X"02",X"DD",X"77",X"01",X"DD",X"7E",X"02",X"E6",
		X"0F",X"FE",X"06",X"38",X"1D",X"47",X"3A",X"58",X"F0",X"FE",X"05",X"38",X"05",X"DD",X"36",X"1F",
		X"0F",X"C9",X"DD",X"7E",X"0C",X"FE",X"80",X"30",X"0A",X"DD",X"7E",X"01",X"EE",X"02",X"DD",X"77",
		X"01",X"C9",X"47",X"3A",X"06",X"F0",X"DD",X"BE",X"09",X"20",X"5E",X"78",X"FE",X"01",X"28",X"1A",
		X"30",X"20",X"21",X"59",X"B9",X"CD",X"EE",X"3D",X"3A",X"8E",X"F3",X"FE",X"02",X"38",X"4A",X"21",
		X"E7",X"F0",X"7E",X"B7",X"20",X"43",X"36",X"80",X"18",X"3F",X"21",X"52",X"B9",X"CD",X"EE",X"3D",
		X"18",X"37",X"3A",X"03",X"F0",X"B7",X"20",X"31",X"3A",X"06",X"F0",X"FE",X"02",X"30",X"2A",X"78",
		X"FE",X"02",X"28",X"25",X"21",X"28",X"F0",X"3A",X"8E",X"F3",X"3C",X"CB",X"27",X"C6",X"08",X"86",
		X"77",X"3A",X"5E",X"F0",X"B7",X"28",X"12",X"AF",X"32",X"5E",X"F0",X"3A",X"5D",X"F0",X"B7",X"20",
		X"08",X"3A",X"12",X"F0",X"EE",X"04",X"32",X"12",X"F0",X"3A",X"15",X"F0",X"B7",X"28",X"0C",X"DD",
		X"36",X"1F",X"0D",X"DD",X"7E",X"04",X"CB",X"2F",X"C3",X"34",X"81",X"3A",X"54",X"F0",X"FE",X"8E",
		X"C2",X"B8",X"80",X"DD",X"36",X"1F",X"01",X"C9",X"DD",X"7E",X"04",X"CB",X"7F",X"3E",X"08",X"28",
		X"02",X"3E",X"EC",X"DD",X"86",X"05",X"4F",X"DD",X"46",X"07",X"CD",X"21",X"72",X"7E",X"FE",X"F0",
		X"28",X"1B",X"FE",X"B0",X"28",X"17",X"FE",X"A9",X"28",X"17",X"FE",X"E9",X"28",X"13",X"FE",X"A2",
		X"28",X"13",X"FE",X"E2",X"28",X"0F",X"DD",X"36",X"1F",X"0A",X"C3",X"0C",X"81",X"0E",X"EF",X"18",
		X"06",X"0E",X"E8",X"18",X"02",X"0E",X"9F",X"DD",X"7E",X"07",X"FE",X"F0",X"30",X"05",X"FE",X"08",
		X"38",X"01",X"71",X"0E",X"12",X"CD",X"4E",X"3D",X"DD",X"36",X"1F",X"01",X"3A",X"06",X"F0",X"DD",
		X"BE",X"09",X"28",X"15",X"3A",X"55",X"F0",X"CB",X"5F",X"20",X"0E",X"E6",X"0F",X"FE",X"06",X"38",
		X"08",X"3E",X"02",X"20",X"0F",X"ED",X"44",X"18",X"0B",X"DD",X"7E",X"04",X"CB",X"7F",X"3E",X"05",
		X"28",X"02",X"ED",X"44",X"DD",X"77",X"04",X"C9",X"DD",X"34",X"1F",X"C3",X"6C",X"83",X"DD",X"34",
		X"1F",X"3A",X"15",X"F0",X"B7",X"20",X"71",X"DD",X"4E",X"05",X"DD",X"46",X"07",X"CD",X"21",X"72",
		X"7E",X"FE",X"EF",X"28",X"0E",X"FE",X"AF",X"28",X"0A",X"FE",X"F0",X"28",X"06",X"FE",X"B0",X"28",
		X"02",X"18",X"55",X"DD",X"36",X"06",X"64",X"DD",X"36",X"1D",X"65",X"DD",X"36",X"16",X"7F",X"DD",
		X"7E",X"07",X"D6",X"10",X"DD",X"77",X"07",X"DD",X"7E",X"02",X"F6",X"10",X"DD",X"77",X"02",X"FD",
		X"21",X"F4",X"F8",X"11",X"04",X"00",X"FD",X"36",X"02",X"66",X"DD",X"46",X"07",X"FD",X"70",X"03",
		X"DD",X"7E",X"05",X"D6",X"10",X"FD",X"77",X"00",X"FD",X"19",X"FD",X"36",X"02",X"67",X"FD",X"77",
		X"00",X"78",X"C6",X"10",X"FD",X"77",X"03",X"DD",X"36",X"03",X"00",X"DD",X"7E",X"01",X"F6",X"01",
		X"DD",X"77",X"01",X"DD",X"36",X"09",X"03",X"C9",X"0E",X"12",X"CD",X"4E",X"3D",X"DD",X"36",X"03",
		X"00",X"DD",X"7E",X"01",X"F6",X"01",X"DD",X"77",X"01",X"DD",X"36",X"1F",X"10",X"C9",X"DD",X"34",
		X"1F",X"FD",X"21",X"F4",X"F8",X"11",X"04",X"00",X"FD",X"36",X"02",X"66",X"DD",X"46",X"07",X"FD",
		X"70",X"03",X"DD",X"7E",X"05",X"D6",X"10",X"FD",X"77",X"00",X"FD",X"19",X"FD",X"36",X"02",X"67",
		X"FD",X"77",X"00",X"78",X"C6",X"10",X"FD",X"77",X"03",X"C9",X"1E",X"00",X"FD",X"21",X"8B",X"F2",
		X"7B",X"FE",X"06",X"CA",X"6C",X"83",X"FD",X"7E",X"00",X"DD",X"BE",X"00",X"CA",X"63",X"83",X"FD",
		X"7E",X"01",X"E6",X"80",X"CA",X"63",X"83",X"FD",X"7E",X"08",X"B7",X"C2",X"63",X"83",X"FD",X"7E",
		X"05",X"B7",X"CA",X"63",X"83",X"47",X"C6",X"0E",X"DD",X"BE",X"05",X"DA",X"63",X"83",X"DD",X"7E",
		X"05",X"C6",X"0E",X"B8",X"DA",X"63",X"83",X"FD",X"7E",X"07",X"47",X"FD",X"86",X"0E",X"38",X"08",
		X"D6",X"04",X"DD",X"BE",X"07",X"DA",X"63",X"83",X"DD",X"7E",X"07",X"DD",X"86",X"0E",X"38",X"06",
		X"D6",X"04",X"B8",X"DA",X"63",X"83",X"0E",X"12",X"CD",X"4E",X"3D",X"3E",X"07",X"DD",X"BE",X"0F",
		X"28",X"0D",X"FD",X"BE",X"0F",X"20",X"68",X"DD",X"E5",X"FD",X"E5",X"DD",X"E1",X"FD",X"E1",X"FD",
		X"BE",X"0F",X"20",X"11",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"06",X"30",X"08",X"DD",X"E5",X"FD",
		X"E5",X"DD",X"E1",X"FD",X"E1",X"DD",X"7E",X"05",X"FD",X"BE",X"05",X"3E",X"02",X"38",X"02",X"ED",
		X"44",X"DD",X"86",X"04",X"FD",X"77",X"04",X"FD",X"7E",X"0C",X"C6",X"04",X"FD",X"77",X"0C",X"FD",
		X"7E",X"07",X"DD",X"BE",X"07",X"30",X"0F",X"D6",X"04",X"FD",X"77",X"07",X"DD",X"7E",X"03",X"C6",
		X"02",X"FD",X"77",X"03",X"18",X"13",X"C6",X"04",X"FD",X"77",X"07",X"FD",X"7E",X"03",X"FE",X"02",
		X"30",X"02",X"3E",X"02",X"D6",X"02",X"FD",X"77",X"03",X"FD",X"36",X"0D",X"08",X"18",X"78",X"DD",
		X"7E",X"05",X"FD",X"BE",X"05",X"30",X"04",X"C6",X"14",X"18",X"02",X"D6",X"14",X"FD",X"77",X"05",
		X"DD",X"7E",X"04",X"FD",X"46",X"04",X"B8",X"20",X"04",X"3C",X"3C",X"05",X"05",X"DD",X"70",X"04",
		X"FD",X"77",X"04",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"28",X"2F",X"CB",X"27",X"47",X"DD",X"86",
		X"07",X"DD",X"77",X"07",X"FD",X"7E",X"07",X"90",X"FD",X"77",X"07",X"DD",X"7E",X"03",X"FE",X"02",
		X"30",X"02",X"3E",X"02",X"D6",X"02",X"47",X"FD",X"7E",X"03",X"FE",X"02",X"30",X"02",X"3E",X"02",
		X"D6",X"02",X"DD",X"77",X"03",X"FD",X"70",X"03",X"18",X"10",X"DD",X"7E",X"07",X"FD",X"BE",X"07",
		X"38",X"05",X"FD",X"34",X"03",X"18",X"03",X"DD",X"34",X"03",X"DD",X"7E",X"0F",X"FD",X"BE",X"0F",
		X"C8",X"30",X"04",X"DD",X"E5",X"FD",X"E1",X"FD",X"7E",X"02",X"FE",X"02",X"C0",X"FD",X"7E",X"01",
		X"47",X"E6",X"0A",X"C0",X"78",X"F6",X"0A",X"FD",X"77",X"01",X"FD",X"36",X"20",X"18",X"FD",X"36",
		X"16",X"00",X"C9",X"01",X"23",X"00",X"FD",X"09",X"1C",X"C3",X"00",X"82",X"01",X"23",X"00",X"DD",
		X"09",X"14",X"7A",X"FE",X"06",X"C2",X"9F",X"7F",X"3A",X"15",X"F0",X"B7",X"C2",X"15",X"84",X"06",
		X"02",X"FD",X"21",X"60",X"F8",X"FD",X"7E",X"00",X"B7",X"28",X"48",X"0E",X"00",X"DD",X"21",X"8B",
		X"F2",X"DD",X"7E",X"01",X"E6",X"80",X"28",X"30",X"DD",X"7E",X"02",X"E6",X"0F",X"28",X"29",X"DD",
		X"7E",X"08",X"B7",X"20",X"23",X"DD",X"7E",X"05",X"D6",X"06",X"FD",X"BE",X"00",X"30",X"19",X"DD",
		X"86",X"0E",X"FD",X"BE",X"00",X"38",X"11",X"DD",X"7E",X"07",X"D6",X"10",X"FD",X"BE",X"03",X"30",
		X"07",X"C6",X"20",X"FD",X"BE",X"03",X"30",X"13",X"11",X"23",X"00",X"DD",X"19",X"0C",X"79",X"FE",
		X"06",X"20",X"BE",X"11",X"04",X"00",X"FD",X"19",X"10",X"AB",X"C9",X"FD",X"36",X"00",X"00",X"FD",
		X"36",X"03",X"00",X"0E",X"37",X"CD",X"4E",X"3D",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"05",X"D0",
		X"DD",X"7E",X"01",X"47",X"E6",X"0A",X"C0",X"78",X"F6",X"0A",X"DD",X"77",X"01",X"DD",X"36",X"16",
		X"7F",X"DD",X"36",X"20",X"18",X"DD",X"7E",X"18",X"B7",X"C8",X"67",X"DD",X"6E",X"17",X"36",X"00",
		X"DD",X"36",X"18",X"00",X"C9",X"3A",X"C2",X"F0",X"B7",X"C8",X"FD",X"21",X"60",X"F8",X"0E",X"02",
		X"21",X"C8",X"F0",X"FD",X"7E",X"00",X"B7",X"28",X"6E",X"7E",X"FE",X"FF",X"28",X"69",X"06",X"06",
		X"DD",X"21",X"8B",X"F2",X"DD",X"7E",X"01",X"E6",X"80",X"28",X"55",X"DD",X"7E",X"08",X"B7",X"20",
		X"4F",X"FD",X"7E",X"00",X"C6",X"08",X"57",X"DD",X"7E",X"05",X"C6",X"08",X"92",X"30",X"02",X"ED",
		X"44",X"FE",X"07",X"30",X"3B",X"FD",X"7E",X"03",X"86",X"57",X"DD",X"7E",X"0E",X"CB",X"3F",X"5F",
		X"DD",X"86",X"07",X"92",X"30",X"02",X"ED",X"44",X"BB",X"30",X"25",X"DD",X"7E",X"01",X"F6",X"03",
		X"DD",X"77",X"01",X"DD",X"36",X"1F",X"10",X"FD",X"36",X"02",X"39",X"36",X"FF",X"23",X"36",X"06",
		X"0E",X"4C",X"3A",X"C2",X"F0",X"FE",X"02",X"DC",X"4E",X"3D",X"0E",X"15",X"CD",X"4E",X"3D",X"C9",
		X"11",X"23",X"00",X"DD",X"19",X"10",X"9D",X"0D",X"C8",X"FD",X"21",X"64",X"F8",X"21",X"CA",X"F0",
		X"18",X"81",X"16",X"00",X"DD",X"21",X"8B",X"F2",X"DD",X"7E",X"01",X"E6",X"81",X"FE",X"81",X"20",
		X"1C",X"DD",X"7E",X"1F",X"D6",X"10",X"38",X"15",X"CD",X"B6",X"88",X"47",X"CB",X"27",X"80",X"21",
		X"2C",X"85",X"85",X"30",X"01",X"24",X"6F",X"E9",X"0E",X"18",X"CD",X"4E",X"3D",X"14",X"7A",X"FE",
		X"06",X"C8",X"01",X"23",X"00",X"DD",X"09",X"18",X"CF",X"DD",X"7E",X"13",X"B7",X"28",X"42",X"67",
		X"DD",X"6E",X"12",X"E5",X"FD",X"E1",X"DD",X"7E",X"07",X"DD",X"86",X"11",X"18",X"13",X"DD",X"7E",
		X"15",X"B7",X"28",X"2D",X"67",X"DD",X"6E",X"14",X"E5",X"FD",X"E1",X"DD",X"7E",X"07",X"DD",X"86",
		X"0A",X"FD",X"77",X"03",X"67",X"DD",X"7E",X"08",X"B7",X"7C",X"28",X"08",X"FE",X"F7",X"30",X"0A",
		X"3E",X"01",X"18",X"09",X"FE",X"F7",X"3E",X"01",X"30",X"03",X"DD",X"7E",X"05",X"FD",X"77",X"00",
		X"C9",X"C1",X"DD",X"36",X"05",X"00",X"DD",X"36",X"03",X"00",X"18",X"A1",X"C3",X"50",X"85",X"C3",
		X"C8",X"85",X"C3",X"21",X"86",X"C3",X"7A",X"86",X"C3",X"B3",X"86",X"C3",X"F6",X"86",X"C3",X"23",
		X"87",X"C3",X"6F",X"87",X"C3",X"DD",X"87",X"C3",X"0C",X"88",X"C3",X"3B",X"88",X"C3",X"76",X"88",
		X"0E",X"00",X"DD",X"7E",X"13",X"B7",X"28",X"0B",X"67",X"DD",X"6E",X"12",X"36",X"00",X"DD",X"36",
		X"13",X"00",X"0C",X"DD",X"7E",X"15",X"B7",X"28",X"0B",X"67",X"DD",X"6E",X"14",X"36",X"00",X"DD",
		X"36",X"15",X"00",X"0C",X"79",X"B7",X"28",X"1B",X"DD",X"7E",X"02",X"4F",X"E6",X"80",X"28",X"08",
		X"79",X"EE",X"80",X"DD",X"77",X"02",X"18",X"0B",X"21",X"51",X"F0",X"35",X"20",X"05",X"0E",X"32",
		X"CD",X"4E",X"3D",X"D5",X"CD",X"EF",X"1B",X"D1",X"DA",X"CD",X"84",X"0E",X"17",X"CD",X"4E",X"3D",
		X"FD",X"E5",X"E1",X"DD",X"75",X"12",X"DD",X"74",X"13",X"DD",X"34",X"1F",X"DD",X"36",X"20",X"04",
		X"3E",X"FD",X"DD",X"77",X"11",X"DD",X"86",X"07",X"FD",X"77",X"03",X"FD",X"36",X"02",X"34",X"DD",
		X"7E",X"05",X"FD",X"77",X"00",X"C3",X"CD",X"84",X"CD",X"D9",X"84",X"DD",X"35",X"20",X"C2",X"CD",
		X"84",X"FD",X"7E",X"02",X"3C",X"FE",X"37",X"30",X"0A",X"FD",X"77",X"02",X"DD",X"36",X"20",X"04",
		X"C3",X"CD",X"84",X"DD",X"36",X"06",X"39",X"3E",X"04",X"2F",X"DD",X"A6",X"01",X"DD",X"77",X"01",
		X"FD",X"7E",X"03",X"C6",X"02",X"FD",X"77",X"03",X"DD",X"36",X"11",X"00",X"DD",X"7E",X"02",X"E6",
		X"10",X"20",X"14",X"DD",X"7E",X"18",X"B7",X"28",X"0A",X"67",X"DD",X"6E",X"17",X"36",X"00",X"DD",
		X"36",X"18",X"00",X"DD",X"36",X"16",X"7F",X"DD",X"36",X"20",X"04",X"DD",X"34",X"1F",X"C3",X"CD",
		X"84",X"CD",X"D9",X"84",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",X"7E",X"02",X"E6",X"10",X"20",
		X"11",X"FD",X"36",X"00",X"00",X"DD",X"34",X"06",X"DD",X"36",X"20",X"04",X"DD",X"34",X"1F",X"C3",
		X"CD",X"84",X"DD",X"36",X"20",X"01",X"D5",X"CD",X"EF",X"1B",X"D1",X"DA",X"CD",X"84",X"FD",X"E5",
		X"E1",X"DD",X"75",X"14",X"DD",X"74",X"15",X"DD",X"34",X"1F",X"DD",X"36",X"20",X"03",X"3E",X"06",
		X"DD",X"77",X"0A",X"DD",X"86",X"07",X"FD",X"77",X"03",X"FD",X"36",X"02",X"37",X"DD",X"7E",X"05",
		X"FD",X"77",X"00",X"DD",X"36",X"06",X"00",X"C3",X"CD",X"84",X"DD",X"7E",X"02",X"E6",X"10",X"20",
		X"18",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",X"36",X"20",X"04",X"DD",X"34",X"06",X"DD",X"7E",
		X"06",X"FE",X"3D",X"D4",X"32",X"3F",X"C3",X"C8",X"84",X"CD",X"D9",X"84",X"CD",X"EE",X"84",X"DD",
		X"35",X"20",X"C2",X"CD",X"84",X"DD",X"36",X"20",X"04",X"DD",X"36",X"0A",X"08",X"DD",X"34",X"1F",
		X"C3",X"CD",X"84",X"CD",X"D9",X"84",X"CD",X"EE",X"84",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",
		X"36",X"20",X"04",X"DD",X"34",X"1F",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"01",X"28",X"04",X"FE",
		X"04",X"20",X"18",X"DD",X"36",X"1D",X"00",X"DD",X"7E",X"18",X"B7",X"28",X"0E",X"67",X"DD",X"6E",
		X"17",X"36",X"00",X"DD",X"36",X"18",X"00",X"DD",X"36",X"16",X"7F",X"DD",X"36",X"11",X"02",X"DD",
		X"36",X"0A",X"0B",X"C3",X"CD",X"84",X"CD",X"D9",X"84",X"CD",X"EE",X"84",X"DD",X"35",X"20",X"C2",
		X"CD",X"84",X"DD",X"36",X"20",X"04",X"DD",X"34",X"1F",X"DD",X"36",X"11",X"04",X"DD",X"7E",X"02",
		X"E6",X"0F",X"FE",X"01",X"CA",X"CD",X"84",X"FE",X"04",X"CA",X"CD",X"84",X"DD",X"36",X"0A",X"0E",
		X"C3",X"CD",X"84",X"CD",X"D9",X"84",X"CD",X"EE",X"84",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",
		X"36",X"20",X"04",X"DD",X"34",X"1F",X"DD",X"7E",X"02",X"E6",X"0F",X"FE",X"01",X"28",X"04",X"FE",
		X"04",X"20",X"21",X"FD",X"36",X"00",X"00",X"DD",X"36",X"0A",X"00",X"DD",X"36",X"11",X"08",X"DD",
		X"7E",X"13",X"B7",X"CA",X"CD",X"84",X"67",X"DD",X"6E",X"12",X"E5",X"FD",X"E1",X"FD",X"36",X"02",
		X"39",X"C3",X"CD",X"84",X"DD",X"36",X"11",X"06",X"DD",X"36",X"0A",X"12",X"C3",X"CD",X"84",X"CD",
		X"D9",X"84",X"DD",X"7E",X"0A",X"B7",X"28",X"43",X"CD",X"EE",X"84",X"DD",X"35",X"20",X"C2",X"CD",
		X"84",X"DD",X"36",X"20",X"04",X"DD",X"34",X"1F",X"DD",X"36",X"1D",X"39",X"DD",X"36",X"11",X"08",
		X"DD",X"7E",X"18",X"B7",X"28",X"0E",X"67",X"DD",X"6E",X"17",X"36",X"00",X"DD",X"36",X"18",X"00",
		X"DD",X"36",X"16",X"7F",X"DD",X"7E",X"02",X"E6",X"0F",X"CA",X"CD",X"84",X"DD",X"36",X"0A",X"14",
		X"FD",X"21",X"68",X"F8",X"FD",X"36",X"00",X"00",X"C3",X"CD",X"84",X"DD",X"35",X"20",X"C2",X"CD",
		X"84",X"FD",X"7E",X"02",X"3C",X"FE",X"3D",X"30",X"0A",X"FD",X"77",X"02",X"DD",X"36",X"20",X"04",
		X"C3",X"CD",X"84",X"AF",X"FD",X"77",X"00",X"CD",X"32",X"3F",X"C3",X"C8",X"84",X"CD",X"D9",X"84",
		X"CD",X"EE",X"84",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",X"36",X"20",X"04",X"DD",X"34",X"1F",
		X"DD",X"36",X"11",X"0A",X"DD",X"7E",X"02",X"E6",X"0F",X"20",X"07",X"DD",X"36",X"0A",X"10",X"C3",
		X"CD",X"84",X"DD",X"34",X"1D",X"DD",X"36",X"0A",X"12",X"C3",X"CD",X"84",X"CD",X"D9",X"84",X"CD",
		X"EE",X"84",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",X"36",X"20",X"04",X"DD",X"34",X"1F",X"DD",
		X"7E",X"02",X"E6",X"0F",X"20",X"0B",X"FD",X"36",X"00",X"00",X"DD",X"36",X"0A",X"00",X"C3",X"CD",
		X"84",X"DD",X"34",X"1D",X"DD",X"36",X"11",X"0C",X"C3",X"CD",X"84",X"CD",X"D9",X"84",X"DD",X"7E",
		X"0A",X"B7",X"28",X"17",X"CD",X"EE",X"84",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",X"36",X"20",
		X"04",X"DD",X"34",X"1F",X"FD",X"36",X"00",X"00",X"C3",X"CD",X"84",X"DD",X"35",X"20",X"C2",X"CD",
		X"84",X"DD",X"36",X"20",X"04",X"DD",X"34",X"1F",X"FD",X"36",X"00",X"00",X"DD",X"36",X"11",X"00",
		X"DD",X"34",X"1D",X"C3",X"CD",X"84",X"DD",X"7E",X"11",X"B7",X"28",X"18",X"CD",X"D9",X"84",X"DD",
		X"35",X"20",X"C2",X"CD",X"84",X"FD",X"36",X"00",X"00",X"DD",X"36",X"11",X"00",X"DD",X"36",X"20",
		X"04",X"C3",X"CD",X"84",X"DD",X"35",X"20",X"C2",X"CD",X"84",X"DD",X"7E",X"1D",X"3C",X"FE",X"3D",
		X"30",X"0A",X"DD",X"77",X"1D",X"DD",X"36",X"20",X"04",X"C3",X"CD",X"84",X"AF",X"FD",X"77",X"00",
		X"CD",X"32",X"3F",X"C3",X"C8",X"84",X"F5",X"D5",X"CD",X"30",X"20",X"38",X"4F",X"DD",X"7E",X"04",
		X"CB",X"7F",X"3E",X"08",X"28",X"02",X"3E",X"EC",X"DD",X"86",X"05",X"4F",X"DD",X"46",X"07",X"CD",
		X"21",X"72",X"7E",X"FE",X"F0",X"28",X"16",X"FE",X"B0",X"28",X"12",X"FE",X"A9",X"28",X"0E",X"FE",
		X"E9",X"28",X"0A",X"FE",X"A2",X"28",X"06",X"FE",X"E2",X"28",X"02",X"18",X"1F",X"0E",X"12",X"CD",
		X"4E",X"3D",X"DD",X"7E",X"04",X"ED",X"44",X"47",X"DD",X"86",X"05",X"DD",X"77",X"05",X"78",X"CB",
		X"2F",X"DD",X"77",X"04",X"DD",X"7E",X"03",X"CB",X"2F",X"DD",X"77",X"03",X"D1",X"F1",X"C9",X"FB",
		X"21",X"A6",X"F0",X"36",X"13",X"21",X"03",X"C9",X"CD",X"07",X"3D",X"DB",X"00",X"E6",X"80",X"CA",
		X"0B",X"A3",X"AF",X"32",X"2A",X"F4",X"F3",X"CD",X"93",X"01",X"FB",X"CD",X"F9",X"3C",X"AF",X"32",
		X"16",X"F4",X"CD",X"B4",X"8B",X"CD",X"3A",X"3D",X"CD",X"25",X"3D",X"CD",X"BE",X"11",X"AF",X"32",
		X"02",X"F4",X"11",X"07",X"B9",X"21",X"F4",X"E9",X"CD",X"18",X"3F",X"11",X"14",X"B9",X"21",X"BB",
		X"EB",X"CD",X"18",X"3F",X"3A",X"2F",X"F4",X"F6",X"30",X"32",X"B2",X"EB",X"E6",X"0F",X"32",X"11",
		X"F4",X"21",X"03",X"F4",X"36",X"80",X"3A",X"2F",X"F4",X"B7",X"C2",X"15",X"8A",X"CD",X"F9",X"3C",
		X"CD",X"DF",X"8B",X"21",X"03",X"F4",X"35",X"20",X"ED",X"3A",X"02",X"F4",X"CB",X"27",X"21",X"E1",
		X"89",X"85",X"30",X"01",X"24",X"6F",X"E9",X"21",X"02",X"F4",X"34",X"CD",X"F9",X"3C",X"CD",X"3A",
		X"3D",X"CD",X"25",X"3D",X"AF",X"32",X"01",X"F4",X"CD",X"BE",X"11",X"F3",X"CD",X"93",X"01",X"FB",
		X"CD",X"F9",X"3C",X"CD",X"B4",X"8B",X"3A",X"2F",X"F4",X"B7",X"CA",X"42",X"89",X"11",X"14",X"B9",
		X"21",X"BB",X"EB",X"CD",X"18",X"3F",X"AF",X"32",X"11",X"F4",X"18",X"59",X"CD",X"F9",X"3C",X"3A",
		X"5E",X"F3",X"B7",X"20",X"12",X"3A",X"2F",X"F4",X"B7",X"28",X"03",X"F1",X"18",X"B9",X"DB",X"00",
		X"E6",X"80",X"C0",X"F1",X"C3",X"0B",X"A3",X"DB",X"01",X"E6",X"04",X"C0",X"F1",X"F1",X"C3",X"26",
		X"89",X"18",X"08",X"18",X"0B",X"18",X"0E",X"18",X"11",X"18",X"14",X"CD",X"5A",X"98",X"18",X"97",
		X"CD",X"54",X"9D",X"18",X"92",X"CD",X"59",X"93",X"18",X"8D",X"CD",X"2E",X"90",X"18",X"88",X"DB",
		X"03",X"E6",X"02",X"20",X"05",X"21",X"A6",X"F0",X"36",X"12",X"21",X"02",X"F4",X"36",X"00",X"23",
		X"36",X"B0",X"C3",X"66",X"89",X"3E",X"01",X"32",X"5D",X"F0",X"3A",X"12",X"F0",X"F6",X"04",X"32",
		X"12",X"F0",X"3E",X"01",X"32",X"6D",X"F3",X"32",X"5E",X"F3",X"21",X"5D",X"F0",X"35",X"20",X"54",
		X"36",X"10",X"3A",X"5C",X"F0",X"EE",X"04",X"32",X"5C",X"F0",X"21",X"5E",X"F3",X"35",X"20",X"44",
		X"36",X"06",X"3A",X"6D",X"F3",X"EE",X"01",X"32",X"6D",X"F3",X"20",X"1D",X"21",X"92",X"E9",X"11",
		X"A9",X"B8",X"CD",X"18",X"3F",X"21",X"F7",X"E9",X"11",X"B2",X"B8",X"CD",X"18",X"3F",X"21",X"57",
		X"EA",X"11",X"C5",X"B8",X"CD",X"18",X"3F",X"18",X"1B",X"21",X"92",X"E9",X"11",X"D8",X"B8",X"CD",
		X"18",X"3F",X"21",X"F7",X"E9",X"11",X"E1",X"B8",X"CD",X"18",X"3F",X"21",X"57",X"EA",X"11",X"F4",
		X"B8",X"CD",X"18",X"3F",X"CD",X"F9",X"3C",X"CD",X"DF",X"8B",X"21",X"11",X"F4",X"3A",X"2F",X"F4",
		X"BE",X"28",X"08",X"32",X"11",X"F4",X"F6",X"30",X"32",X"B2",X"EB",X"DB",X"01",X"2F",X"E6",X"04",
		X"20",X"33",X"3A",X"7E",X"F0",X"FE",X"04",X"38",X"81",X"3A",X"5C",X"F0",X"F6",X"04",X"32",X"5C",
		X"F0",X"21",X"C5",X"8A",X"E5",X"3A",X"2A",X"F4",X"6F",X"CB",X"27",X"85",X"21",X"CC",X"8A",X"85",
		X"30",X"01",X"24",X"6F",X"E9",X"21",X"2A",X"F4",X"34",X"C3",X"26",X"89",X"C3",X"59",X"93",X"C3",
		X"35",X"94",X"C3",X"9D",X"97",X"AF",X"32",X"2A",X"F4",X"CD",X"F9",X"3C",X"CD",X"DF",X"8B",X"3A",
		X"2F",X"F4",X"3D",X"32",X"2F",X"F4",X"F6",X"30",X"32",X"B2",X"EB",X"CD",X"F9",X"3C",X"CD",X"DF",
		X"8B",X"AF",X"32",X"5D",X"F0",X"3A",X"12",X"F0",X"EE",X"04",X"32",X"12",X"F0",X"21",X"A6",X"F0",
		X"36",X"12",X"06",X"E0",X"21",X"81",X"E9",X"36",X"00",X"23",X"10",X"FB",X"CD",X"F9",X"3C",X"CD",
		X"DF",X"8B",X"21",X"03",X"F0",X"36",X"01",X"21",X"B0",X"F0",X"36",X"02",X"21",X"35",X"F0",X"36",
		X"00",X"CD",X"F9",X"3C",X"CD",X"DF",X"8B",X"3E",X"09",X"06",X"03",X"21",X"7F",X"F3",X"77",X"23",
		X"10",X"FC",X"F6",X"30",X"06",X"03",X"21",X"6E",X"E8",X"77",X"23",X"10",X"FC",X"AF",X"06",X"0A",
		X"21",X"B2",X"EB",X"77",X"23",X"10",X"FC",X"0E",X"02",X"CD",X"4E",X"3D",X"AF",X"32",X"2E",X"F0",
		X"CD",X"F9",X"3C",X"CD",X"DF",X"8B",X"3A",X"03",X"F0",X"47",X"E6",X"80",X"20",X"37",X"78",X"B7",
		X"20",X"EA",X"3A",X"7A",X"F3",X"B7",X"20",X"E4",X"3A",X"06",X"F0",X"FE",X"02",X"30",X"0C",X"3A",
		X"09",X"F0",X"B7",X"20",X"06",X"3A",X"82",X"F0",X"B7",X"20",X"D1",X"3A",X"2E",X"F0",X"FE",X"80",
		X"38",X"0D",X"3A",X"43",X"F0",X"B7",X"20",X"C8",X"3E",X"02",X"32",X"43",X"F0",X"18",X"BD",X"3C",
		X"32",X"2E",X"F0",X"18",X"BB",X"CD",X"19",X"8C",X"3A",X"2F",X"F4",X"B7",X"CA",X"3E",X"89",X"11",
		X"14",X"B9",X"21",X"BB",X"EB",X"CD",X"18",X"3F",X"AF",X"32",X"11",X"F4",X"0E",X"02",X"CD",X"4E",
		X"3D",X"C3",X"15",X"8A",X"C5",X"0E",X"30",X"3A",X"14",X"F0",X"B7",X"28",X"02",X"0E",X"0D",X"11",
		X"41",X"B9",X"21",X"47",X"E8",X"CD",X"18",X"3F",X"06",X"06",X"21",X"6A",X"E8",X"11",X"39",X"F4",
		X"1A",X"B7",X"28",X"01",X"81",X"77",X"2B",X"13",X"1A",X"81",X"77",X"10",X"F9",X"C1",X"C9",X"CD",
		X"B9",X"2A",X"CD",X"40",X"1C",X"CD",X"A6",X"4B",X"CD",X"96",X"72",X"CD",X"CC",X"27",X"CD",X"B5",
		X"79",X"CD",X"99",X"7F",X"CD",X"34",X"32",X"CD",X"A2",X"84",X"CD",X"40",X"4C",X"CD",X"A0",X"52",
		X"CD",X"1D",X"54",X"CD",X"7E",X"5E",X"CD",X"1E",X"5A",X"CD",X"4F",X"23",X"CD",X"15",X"24",X"CD",
		X"85",X"55",X"CD",X"1E",X"63",X"CD",X"52",X"64",X"C9",X"CD",X"F9",X"3C",X"F3",X"CD",X"93",X"01",
		X"FB",X"21",X"F3",X"E9",X"11",X"1C",X"B9",X"CD",X"18",X"3F",X"21",X"05",X"F4",X"36",X"80",X"06",
		X"07",X"21",X"82",X"F3",X"11",X"39",X"F4",X"1A",X"BE",X"38",X"08",X"20",X"14",X"13",X"23",X"10",
		X"F6",X"18",X"0E",X"21",X"82",X"F3",X"11",X"39",X"F4",X"06",X"07",X"7E",X"12",X"23",X"13",X"10",
		X"FA",X"CD",X"B4",X"8B",X"CD",X"F9",X"3C",X"CD",X"DF",X"8B",X"21",X"05",X"F4",X"35",X"20",X"F4",
		X"CD",X"3A",X"3D",X"CD",X"F9",X"3C",X"21",X"5D",X"F3",X"CD",X"2E",X"3D",X"CD",X"F9",X"3C",X"21",
		X"F3",X"E9",X"CD",X"15",X"3F",X"CD",X"BE",X"11",X"CD",X"B4",X"8B",X"CD",X"AE",X"A0",X"CD",X"39",
		X"A2",X"CD",X"99",X"A1",X"06",X"78",X"CD",X"F9",X"3C",X"10",X"FB",X"21",X"5D",X"F3",X"36",X"01",
		X"F3",X"CD",X"93",X"01",X"FB",X"3A",X"60",X"F3",X"FE",X"0B",X"30",X"0A",X"CD",X"3C",X"8D",X"06",
		X"1E",X"CD",X"F9",X"3C",X"10",X"FB",X"3A",X"2F",X"F4",X"B7",X"CC",X"2E",X"90",X"F3",X"CD",X"93",
		X"01",X"FB",X"CD",X"F9",X"3C",X"CD",X"B4",X"8B",X"CD",X"F9",X"3C",X"CD",X"3A",X"3D",X"CD",X"25",
		X"3D",X"CD",X"BE",X"11",X"CD",X"F9",X"3C",X"C9",X"55",X"53",X"45",X"20",X"53",X"54",X"45",X"45",
		X"52",X"49",X"4E",X"47",X"20",X"57",X"48",X"45",X"45",X"4C",X"00",X"54",X"4F",X"20",X"53",X"45",
		X"4C",X"45",X"43",X"54",X"20",X"49",X"4E",X"49",X"54",X"49",X"41",X"4C",X"20",X"00",X"55",X"53",
		X"45",X"20",X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"20",X"54",X"52",X"49",X"47",X"47",X"45",
		X"52",X"00",X"54",X"4F",X"20",X"45",X"4E",X"54",X"45",X"52",X"20",X"53",X"45",X"4C",X"45",X"43",
		X"54",X"49",X"4F",X"4E",X"00",X"20",X"45",X"4E",X"54",X"45",X"52",X"20",X"33",X"20",X"49",X"4E",
		X"49",X"54",X"49",X"41",X"4C",X"53",X"20",X"00",X"20",X"43",X"4F",X"4E",X"47",X"52",X"41",X"54",
		X"55",X"4C",X"41",X"54",X"49",X"4F",X"4E",X"53",X"21",X"20",X"20",X"00",X"F3",X"CD",X"93",X"01",
		X"FB",X"CD",X"F9",X"3C",X"21",X"FE",X"F0",X"36",X"FF",X"21",X"E8",X"F0",X"36",X"01",X"21",X"E4",
		X"F0",X"36",X"60",X"21",X"E2",X"F0",X"36",X"76",X"21",X"90",X"E9",X"22",X"9B",X"F0",X"3E",X"41",
		X"06",X"1A",X"21",X"BB",X"EA",X"77",X"3C",X"FE",X"4F",X"20",X"03",X"21",X"5D",X"EB",X"2B",X"2B",
		X"10",X"F3",X"CD",X"E7",X"8F",X"2B",X"2B",X"CD",X"F7",X"8F",X"21",X"97",X"E8",X"11",X"C8",X"8C",
		X"CD",X"18",X"3F",X"21",X"D7",X"E8",X"11",X"DB",X"8C",X"CD",X"18",X"3F",X"21",X"37",X"E9",X"11",
		X"EE",X"8C",X"CD",X"18",X"3F",X"21",X"77",X"E9",X"11",X"02",X"8D",X"CD",X"18",X"3F",X"AF",X"32",
		X"68",X"F3",X"32",X"69",X"F3",X"32",X"6B",X"F3",X"3E",X"08",X"32",X"6A",X"F3",X"DD",X"21",X"FF",
		X"F0",X"21",X"5E",X"F3",X"36",X"FF",X"23",X"36",X"07",X"0E",X"02",X"CD",X"4E",X"3D",X"3A",X"12",
		X"F0",X"F6",X"80",X"32",X"12",X"F0",X"21",X"6D",X"F3",X"36",X"01",X"21",X"6C",X"F3",X"36",X"01",
		X"3A",X"6D",X"F3",X"B7",X"28",X"02",X"18",X"25",X"3A",X"6C",X"F3",X"B7",X"28",X"1F",X"21",X"97",
		X"E8",X"11",X"15",X"8D",X"CD",X"18",X"3F",X"21",X"D7",X"E8",X"CD",X"15",X"3F",X"21",X"37",X"E9",
		X"CD",X"15",X"3F",X"21",X"77",X"E9",X"CD",X"15",X"3F",X"AF",X"32",X"6C",X"F3",X"DB",X"01",X"2F",
		X"E6",X"04",X"C2",X"15",X"8F",X"3A",X"6A",X"F3",X"B7",X"C2",X"DD",X"8E",X"0E",X"00",X"3A",X"A1",
		X"F0",X"47",X"CB",X"7F",X"28",X"02",X"ED",X"44",X"FE",X"03",X"38",X"27",X"D6",X"01",X"4F",X"3A",
		X"69",X"F3",X"B7",X"20",X"1E",X"DD",X"7E",X"00",X"B7",X"20",X"18",X"CB",X"78",X"3A",X"68",X"F3",
		X"20",X"08",X"D6",X"01",X"30",X"0A",X"3E",X"1B",X"18",X"06",X"3C",X"FE",X"1C",X"38",X"01",X"AF",
		X"32",X"68",X"F3",X"3A",X"68",X"F3",X"FE",X"0E",X"21",X"BB",X"EA",X"16",X"B4",X"38",X"07",X"21",
		X"5B",X"EB",X"16",X"DC",X"D6",X"0E",X"5F",X"B7",X"28",X"09",X"CB",X"27",X"ED",X"44",X"85",X"38",
		X"01",X"25",X"6F",X"3A",X"68",X"F3",X"FE",X"1A",X"38",X"1A",X"28",X"0C",X"3A",X"69",X"F3",X"B7",
		X"CC",X"D7",X"8F",X"C4",X"F7",X"8F",X"18",X"2B",X"3A",X"69",X"F3",X"B7",X"CC",X"D7",X"8F",X"C4",
		X"E7",X"8F",X"18",X"1F",X"3A",X"69",X"F3",X"B7",X"28",X"05",X"3A",X"68",X"F3",X"C6",X"41",X"77",
		X"B7",X"28",X"10",X"3A",X"6B",X"F3",X"FE",X"02",X"20",X"09",X"3D",X"32",X"6B",X"F3",X"21",X"68",
		X"F3",X"36",X"1B",X"21",X"01",X"F0",X"72",X"7B",X"CB",X"27",X"CB",X"27",X"CB",X"27",X"CB",X"27",
		X"C6",X"1D",X"32",X"00",X"F0",X"DD",X"21",X"6C",X"F8",X"DD",X"77",X"00",X"DD",X"77",X"04",X"DD",
		X"36",X"02",X"21",X"DD",X"36",X"06",X"22",X"7E",X"DD",X"77",X"03",X"C6",X"10",X"DD",X"77",X"07",
		X"3A",X"69",X"F3",X"EE",X"01",X"32",X"69",X"F3",X"3E",X"08",X"91",X"18",X"01",X"3D",X"32",X"6A",
		X"F3",X"CD",X"F9",X"3C",X"CD",X"40",X"4C",X"3A",X"E8",X"F0",X"B7",X"28",X"21",X"21",X"5E",X"F3",
		X"35",X"C2",X"D0",X"8D",X"23",X"35",X"28",X"06",X"2B",X"36",X"FF",X"C3",X"D0",X"8D",X"3A",X"FF",
		X"F0",X"B7",X"28",X"07",X"34",X"2B",X"36",X"20",X"C3",X"D0",X"8D",X"32",X"E8",X"F0",X"3A",X"69",
		X"F3",X"B7",X"C2",X"D0",X"8D",X"3A",X"12",X"F0",X"EE",X"80",X"32",X"12",X"F0",X"11",X"61",X"F3",
		X"21",X"90",X"E9",X"06",X"03",X"7E",X"12",X"2B",X"2B",X"13",X"10",X"F9",X"AF",X"32",X"6A",X"F3",
		X"32",X"69",X"F3",X"21",X"E4",X"F0",X"36",X"F8",X"21",X"97",X"E8",X"CD",X"15",X"3F",X"21",X"D7",
		X"E8",X"CD",X"15",X"3F",X"21",X"37",X"E9",X"11",X"28",X"8D",X"CD",X"18",X"3F",X"21",X"77",X"E9",
		X"CD",X"15",X"3F",X"DB",X"01",X"2F",X"E6",X"04",X"20",X"6D",X"DD",X"21",X"6C",X"F8",X"0E",X"BC",
		X"16",X"CF",X"1E",X"00",X"CD",X"8E",X"3D",X"3A",X"6A",X"F3",X"B7",X"20",X"14",X"3A",X"69",X"F3",
		X"B7",X"CC",X"07",X"90",X"C4",X"18",X"90",X"3A",X"69",X"F3",X"EE",X"01",X"32",X"69",X"F3",X"3E",
		X"05",X"3D",X"32",X"6A",X"F3",X"21",X"00",X"F0",X"7E",X"FE",X"85",X"28",X"08",X"3E",X"02",X"38",
		X"02",X"ED",X"44",X"86",X"77",X"3A",X"01",X"F0",X"D6",X"02",X"32",X"01",X"F0",X"21",X"E4",X"F0",
		X"BE",X"20",X"0B",X"7E",X"FE",X"F0",X"28",X"1F",X"36",X"F0",X"DD",X"36",X"02",X"00",X"3A",X"00",
		X"F0",X"DD",X"77",X"00",X"DD",X"77",X"04",X"3A",X"01",X"F0",X"DD",X"77",X"03",X"C6",X"10",X"DD",
		X"77",X"07",X"CD",X"F9",X"3C",X"18",X"A0",X"CD",X"6E",X"A0",X"06",X"20",X"CD",X"F9",X"3C",X"10",
		X"FB",X"0E",X"01",X"CD",X"4E",X"3D",X"C9",X"E5",X"FD",X"E1",X"FD",X"36",X"00",X"00",X"FD",X"36",
		X"E0",X"00",X"FD",X"36",X"C0",X"00",X"C9",X"E5",X"FD",X"E1",X"FD",X"36",X"C0",X"52",X"FD",X"36",
		X"E0",X"55",X"FD",X"36",X"00",X"42",X"C9",X"E5",X"FD",X"E1",X"FD",X"36",X"C0",X"45",X"FD",X"36",
		X"E0",X"4E",X"FD",X"36",X"00",X"44",X"C9",X"FD",X"21",X"90",X"E9",X"FD",X"36",X"00",X"00",X"FD",
		X"36",X"FE",X"00",X"FD",X"36",X"FC",X"00",X"C9",X"FD",X"21",X"90",X"E9",X"21",X"61",X"F3",X"7E",
		X"FD",X"77",X"00",X"23",X"7E",X"FD",X"77",X"FE",X"23",X"7E",X"FD",X"77",X"FC",X"C9",X"CD",X"BC",
		X"89",X"21",X"5D",X"F3",X"CD",X"2E",X"3D",X"21",X"5D",X"F3",X"36",X"01",X"F3",X"CD",X"93",X"01",
		X"FB",X"CD",X"3A",X"3D",X"AF",X"32",X"6C",X"F3",X"CD",X"BC",X"89",X"3A",X"6C",X"F3",X"47",X"CB",
		X"27",X"80",X"21",X"6E",X"90",X"85",X"30",X"01",X"24",X"6F",X"E9",X"21",X"6C",X"F3",X"34",X"CD",
		X"ED",X"36",X"CD",X"1E",X"63",X"CD",X"1E",X"5A",X"CD",X"BC",X"89",X"C3",X"4B",X"90",X"C3",X"8C",
		X"90",X"C3",X"AA",X"90",X"C3",X"C3",X"90",X"C3",X"DD",X"90",X"C3",X"00",X"91",X"C3",X"45",X"91",
		X"C3",X"96",X"91",X"C3",X"C6",X"91",X"C3",X"DE",X"91",X"C3",X"FB",X"91",X"21",X"D9",X"F0",X"36",
		X"01",X"21",X"DB",X"F0",X"36",X"03",X"21",X"E2",X"F0",X"36",X"26",X"21",X"E4",X"F0",X"36",X"00",
		X"3A",X"2F",X"F4",X"B7",X"CA",X"5B",X"90",X"C3",X"5B",X"90",X"3A",X"E4",X"F0",X"C6",X"02",X"32",
		X"E4",X"F0",X"FE",X"24",X"DA",X"5F",X"90",X"21",X"93",X"E8",X"11",X"79",X"92",X"CD",X"18",X"3F",
		X"C3",X"5B",X"90",X"3A",X"E4",X"F0",X"C6",X"02",X"32",X"E4",X"F0",X"FE",X"3C",X"DA",X"5F",X"90",
		X"21",X"EE",X"F0",X"36",X"01",X"21",X"00",X"F0",X"36",X"36",X"C3",X"5B",X"90",X"21",X"EE",X"F0",
		X"3A",X"EF",X"F0",X"B6",X"C2",X"5F",X"90",X"DD",X"21",X"40",X"F4",X"FD",X"21",X"F4",X"E8",X"CD",
		X"37",X"92",X"DD",X"21",X"6A",X"F4",X"FD",X"21",X"EF",X"E8",X"CD",X"46",X"92",X"C3",X"5B",X"90",
		X"3A",X"E4",X"F0",X"C6",X"02",X"32",X"E4",X"F0",X"FE",X"5C",X"DA",X"5F",X"90",X"3E",X"5E",X"32",
		X"E4",X"F0",X"21",X"77",X"E9",X"11",X"84",X"92",X"CD",X"18",X"3F",X"21",X"6F",X"F3",X"36",X"7E",
		X"DD",X"21",X"B4",X"E9",X"DD",X"22",X"70",X"F3",X"21",X"6E",X"F3",X"36",X"32",X"DD",X"21",X"43",
		X"F4",X"DD",X"22",X"74",X"F3",X"DD",X"21",X"6E",X"F4",X"DD",X"22",X"72",X"F3",X"21",X"6D",X"F3",
		X"36",X"08",X"C3",X"5B",X"90",X"3A",X"E4",X"F0",X"C6",X"02",X"32",X"E4",X"F0",X"21",X"6F",X"F3",
		X"BE",X"DA",X"5F",X"90",X"C6",X"10",X"77",X"FD",X"2A",X"70",X"F3",X"3A",X"6E",X"F3",X"FD",X"77",
		X"02",X"3C",X"32",X"6E",X"F3",X"DD",X"2A",X"74",X"F3",X"CD",X"37",X"92",X"DD",X"22",X"74",X"F3",
		X"FD",X"2B",X"FD",X"2B",X"DD",X"2A",X"72",X"F3",X"CD",X"46",X"92",X"DD",X"22",X"72",X"F3",X"FD",
		X"2A",X"70",X"F3",X"11",X"40",X"00",X"FD",X"19",X"FD",X"22",X"70",X"F3",X"21",X"6D",X"F3",X"35",
		X"C2",X"5F",X"90",X"C3",X"5B",X"90",X"3A",X"E4",X"F0",X"C6",X"02",X"32",X"E4",X"F0",X"21",X"6F",
		X"F3",X"BE",X"DA",X"5F",X"90",X"FD",X"2A",X"70",X"F3",X"FD",X"36",X"03",X"31",X"FD",X"36",X"02",
		X"30",X"DD",X"2A",X"74",X"F3",X"CD",X"37",X"92",X"FD",X"2B",X"FD",X"2B",X"DD",X"2A",X"72",X"F3",
		X"CD",X"46",X"92",X"C3",X"5B",X"90",X"3A",X"DB",X"F0",X"3C",X"32",X"DB",X"F0",X"FE",X"09",X"CA",
		X"5B",X"90",X"CD",X"BC",X"89",X"CD",X"BC",X"89",X"CD",X"BC",X"89",X"C3",X"5F",X"90",X"3A",X"E4",
		X"F0",X"D6",X"02",X"32",X"E4",X"F0",X"FE",X"02",X"D2",X"5F",X"90",X"3E",X"01",X"32",X"E3",X"F0",
		X"32",X"E1",X"F0",X"21",X"6D",X"F3",X"36",X"F0",X"C3",X"5B",X"90",X"21",X"6D",X"F3",X"35",X"C2",
		X"5F",X"90",X"F3",X"CD",X"93",X"01",X"FB",X"CD",X"F9",X"3C",X"11",X"41",X"B9",X"21",X"47",X"E8",
		X"CD",X"18",X"3F",X"06",X"06",X"21",X"6A",X"E8",X"11",X"39",X"F4",X"1A",X"B7",X"28",X"02",X"F6",
		X"30",X"77",X"2B",X"13",X"1A",X"F6",X"30",X"77",X"10",X"F8",X"CD",X"F9",X"3C",X"CD",X"3A",X"3D",
		X"CD",X"25",X"3D",X"CD",X"BE",X"11",X"C9",X"06",X"03",X"DD",X"7E",X"00",X"FD",X"77",X"00",X"DD",
		X"23",X"FD",X"2B",X"10",X"F4",X"C9",X"DD",X"7E",X"00",X"B7",X"28",X"02",X"F6",X"30",X"FD",X"77",
		X"00",X"06",X"03",X"DD",X"23",X"FD",X"2B",X"DD",X"7E",X"00",X"4F",X"E6",X"F0",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"F6",X"30",X"FD",X"77",X"00",X"79",X"E6",X"0F",X"F6",X"30",X"FD",
		X"77",X"FF",X"FD",X"2B",X"10",X"DD",X"DD",X"23",X"C9",X"54",X"4F",X"50",X"20",X"20",X"41",X"47",
		X"45",X"4E",X"54",X"00",X"53",X"50",X"45",X"43",X"49",X"41",X"4C",X"20",X"46",X"4F",X"52",X"43",
		X"45",X"20",X"54",X"45",X"41",X"4D",X"00",X"20",X"20",X"31",X"53",X"54",X"20",X"53",X"54",X"41",
		X"47",X"45",X"20",X"4F",X"46",X"20",X"47",X"41",X"4D",X"45",X"00",X"20",X"20",X"20",X"52",X"55",
		X"4E",X"53",X"20",X"4F",X"4E",X"20",X"41",X"20",X"54",X"49",X"4D",X"45",X"52",X"00",X"20",X"57",
		X"49",X"54",X"48",X"20",X"55",X"4E",X"4C",X"49",X"4D",X"49",X"54",X"45",X"44",X"20",X"43",X"41",
		X"52",X"53",X"00",X"20",X"41",X"46",X"54",X"45",X"52",X"20",X"54",X"49",X"4D",X"45",X"52",X"20",
		X"45",X"58",X"50",X"49",X"52",X"45",X"53",X"00",X"42",X"41",X"53",X"45",X"53",X"20",X"57",X"49",
		X"4C",X"4C",X"20",X"42",X"45",X"20",X"41",X"57",X"41",X"52",X"44",X"45",X"44",X"00",X"20",X"20",
		X"46",X"4F",X"52",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"20",X"45",X"41",X"52",X"4E",X"45",
		X"44",X"00",X"20",X"20",X"41",X"44",X"44",X"49",X"54",X"49",X"4F",X"4E",X"41",X"4C",X"20",X"42",
		X"41",X"53",X"45",X"53",X"00",X"20",X"57",X"49",X"4C",X"4C",X"20",X"42",X"45",X"20",X"41",X"57",
		X"41",X"52",X"44",X"45",X"44",X"20",X"41",X"54",X"00",X"20",X"20",X"20",X"20",X"20",X"30",X"30",
		X"30",X"20",X"20",X"20",X"20",X"20",X"20",X"30",X"30",X"30",X"00",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"CD",X"3A",X"3D",X"CD",X"BC",X"89",X"21",
		X"5D",X"F3",X"36",X"01",X"F3",X"CD",X"93",X"01",X"FB",X"21",X"98",X"E8",X"11",X"97",X"92",X"CD",
		X"18",X"3F",X"21",X"D8",X"E8",X"11",X"AB",X"92",X"CD",X"18",X"3F",X"21",X"18",X"E9",X"11",X"BE",
		X"92",X"CD",X"18",X"3F",X"21",X"78",X"E9",X"11",X"D3",X"92",X"CD",X"18",X"3F",X"21",X"B8",X"E9",
		X"11",X"E8",X"92",X"CD",X"18",X"3F",X"21",X"F8",X"E9",X"11",X"FE",X"92",X"CD",X"18",X"3F",X"21",
		X"58",X"EA",X"11",X"12",X"93",X"CD",X"18",X"3F",X"21",X"98",X"EA",X"11",X"25",X"93",X"CD",X"18",
		X"3F",X"21",X"D8",X"EA",X"11",X"39",X"93",X"CD",X"18",X"3F",X"21",X"18",X"EB",X"11",X"39",X"93",
		X"CD",X"18",X"3F",X"21",X"58",X"EB",X"11",X"4B",X"93",X"CD",X"18",X"3F",X"21",X"D4",X"EA",X"CD",
		X"EF",X"93",X"CD",X"62",X"3E",X"21",X"CB",X"EA",X"CD",X"EF",X"93",X"CD",X"62",X"3E",X"21",X"14",
		X"EB",X"CD",X"EF",X"93",X"CD",X"62",X"3E",X"21",X"0B",X"EB",X"CD",X"EF",X"93",X"18",X"16",X"11",
		X"7F",X"F2",X"1A",X"F6",X"30",X"77",X"23",X"1B",X"1A",X"F6",X"30",X"77",X"1B",X"1A",X"B7",X"C8",
		X"23",X"F6",X"30",X"77",X"C9",X"06",X"FF",X"CD",X"BC",X"89",X"10",X"FB",X"C9",X"42",X"45",X"57",
		X"41",X"52",X"45",X"20",X"4F",X"46",X"20",X"00",X"42",X"41",X"52",X"52",X"45",X"4C",X"20",X"44",
		X"55",X"4D",X"50",X"45",X"52",X"00",X"44",X"4F",X"43",X"54",X"4F",X"52",X"20",X"54",X"4F",X"52",
		X"50",X"45",X"44",X"4F",X"00",X"CD",X"3A",X"3D",X"CD",X"BC",X"89",X"21",X"5D",X"F3",X"36",X"01",
		X"F3",X"CD",X"93",X"01",X"FB",X"3E",X"04",X"06",X"50",X"21",X"70",X"E3",X"77",X"23",X"10",X"FC",
		X"3E",X"EF",X"06",X"40",X"77",X"23",X"10",X"FC",X"21",X"5B",X"E8",X"11",X"0D",X"94",X"CD",X"18",
		X"3F",X"21",X"51",X"E8",X"11",X"2C",X"9C",X"CD",X"18",X"3F",X"21",X"B9",X"E8",X"11",X"3D",X"9C",
		X"CD",X"18",X"3F",X"21",X"CB",X"E8",X"11",X"33",X"9D",X"CD",X"18",X"3F",X"21",X"39",X"E9",X"11",
		X"62",X"9C",X"CD",X"18",X"3F",X"21",X"4B",X"E9",X"11",X"33",X"9D",X"CD",X"18",X"3F",X"21",X"B9",
		X"E9",X"11",X"86",X"9C",X"CD",X"18",X"3F",X"21",X"CB",X"E9",X"11",X"3E",X"9D",X"CD",X"18",X"3F",
		X"21",X"78",X"EA",X"11",X"AA",X"9C",X"CD",X"18",X"3F",X"21",X"8B",X"EA",X"11",X"49",X"9D",X"CD",
		X"18",X"3F",X"21",X"17",X"EB",X"11",X"18",X"94",X"CD",X"18",X"3F",X"21",X"2B",X"EB",X"11",X"33",
		X"9D",X"CD",X"18",X"3F",X"21",X"97",X"EB",X"11",X"26",X"94",X"CD",X"18",X"3F",X"21",X"AB",X"EB",
		X"11",X"3E",X"9D",X"CD",X"18",X"3F",X"11",X"04",X"00",X"DD",X"21",X"04",X"F8",X"DD",X"36",X"00",
		X"1B",X"DD",X"36",X"01",X"20",X"DD",X"36",X"02",X"0D",X"DD",X"36",X"03",X"42",X"DD",X"19",X"DD",
		X"36",X"00",X"32",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"0D",X"DD",X"36",X"03",X"42",X"DD",
		X"19",X"DD",X"36",X"00",X"23",X"DD",X"36",X"01",X"20",X"DD",X"36",X"02",X"AF",X"DD",X"36",X"03",
		X"C7",X"DD",X"19",X"DD",X"36",X"00",X"29",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"AF",X"DD",
		X"36",X"03",X"C7",X"DD",X"19",X"DD",X"36",X"00",X"22",X"DD",X"36",X"01",X"20",X"DD",X"36",X"02",
		X"AF",X"DD",X"36",X"03",X"E9",X"DD",X"19",X"DD",X"36",X"00",X"2A",X"DD",X"36",X"01",X"00",X"DD",
		X"36",X"02",X"AF",X"DD",X"36",X"03",X"E9",X"DD",X"19",X"DD",X"36",X"00",X"28",X"DD",X"36",X"01",
		X"00",X"DD",X"36",X"02",X"7C",X"DD",X"36",X"03",X"22",X"DD",X"19",X"DD",X"36",X"00",X"28",X"DD",
		X"36",X"01",X"00",X"DD",X"36",X"02",X"7D",X"DD",X"36",X"03",X"32",X"DD",X"19",X"DD",X"36",X"00",
		X"26",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"27",X"DD",X"36",X"03",X"40",X"DD",X"19",X"DD",
		X"36",X"00",X"26",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"28",X"DD",X"36",X"03",X"50",X"DD",
		X"19",X"DD",X"36",X"00",X"26",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"25",X"DD",X"36",X"03",
		X"60",X"DD",X"19",X"DD",X"36",X"00",X"26",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"26",X"DD",
		X"36",X"03",X"70",X"DD",X"19",X"DD",X"36",X"00",X"32",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",
		X"10",X"DD",X"36",X"03",X"70",X"DD",X"19",X"DD",X"36",X"00",X"26",X"DD",X"36",X"01",X"00",X"DD",
		X"36",X"02",X"70",X"DD",X"36",X"03",X"BA",X"DD",X"19",X"DD",X"36",X"00",X"26",X"DD",X"36",X"01",
		X"00",X"DD",X"36",X"02",X"71",X"DD",X"36",X"03",X"CA",X"DD",X"19",X"DD",X"36",X"00",X"27",X"DD",
		X"36",X"01",X"00",X"DD",X"36",X"02",X"74",X"DD",X"36",X"03",X"C1",X"DD",X"19",X"DD",X"36",X"00",
		X"26",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"AB",X"DD",X"36",X"03",X"D8",X"DD",X"19",X"DD",
		X"36",X"00",X"26",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"AC",X"DD",X"36",X"03",X"E8",X"DD",
		X"19",X"DD",X"36",X"00",X"26",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"AD",X"DD",X"36",X"03",
		X"DF",X"DD",X"21",X"D8",X"F9",X"DD",X"36",X"00",X"2E",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",
		X"02",X"DD",X"36",X"03",X"8D",X"3E",X"02",X"32",X"D9",X"F0",X"AF",X"32",X"E3",X"F0",X"32",X"E1",
		X"F0",X"3E",X"09",X"32",X"DB",X"F0",X"3E",X"1E",X"32",X"E2",X"F0",X"3E",X"98",X"32",X"E4",X"F0",
		X"21",X"03",X"F4",X"36",X"04",X"0E",X"02",X"06",X"FF",X"C5",X"CD",X"BC",X"89",X"CD",X"1E",X"5A",
		X"DD",X"21",X"04",X"F8",X"01",X"04",X"00",X"DD",X"7E",X"01",X"EE",X"10",X"DD",X"77",X"01",X"DD",
		X"09",X"DD",X"7E",X"01",X"EE",X"10",X"DD",X"77",X"01",X"21",X"03",X"F4",X"35",X"20",X"1F",X"36",
		X"04",X"DD",X"09",X"3E",X"AF",X"DD",X"BE",X"02",X"20",X"02",X"3E",X"B3",X"DD",X"77",X"02",X"DD",
		X"09",X"DD",X"77",X"02",X"DD",X"09",X"DD",X"77",X"02",X"DD",X"09",X"DD",X"77",X"02",X"C1",X"10",
		X"B8",X"0D",X"20",X"B3",X"C9",X"57",X"45",X"41",X"50",X"4F",X"4E",X"53",X"00",X"4D",X"41",X"59",
		X"20",X"42",X"45",X"20",X"45",X"41",X"52",X"4E",X"45",X"44",X"20",X"42",X"59",X"20",X"45",X"4E",
		X"54",X"45",X"52",X"49",X"4E",X"47",X"00",X"57",X"45",X"41",X"50",X"4F",X"4E",X"53",X"20",X"56",
		X"41",X"4E",X"20",X"57",X"49",X"54",X"48",X"20",X"52",X"41",X"4D",X"50",X"00",X"57",X"45",X"41",
		X"50",X"4F",X"4E",X"53",X"20",X"41",X"56",X"41",X"49",X"4C",X"41",X"42",X"4C",X"45",X"00",X"41",
		X"52",X"45",X"20",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"45",X"44",X"20",X"4F",X"4E",X"20",
		X"43",X"4F",X"4E",X"53",X"4F",X"4C",X"45",X"00",X"57",X"45",X"41",X"50",X"4F",X"4E",X"20",X"53",
		X"45",X"4C",X"45",X"43",X"54",X"49",X"4F",X"4E",X"00",X"4C",X"45",X"46",X"54",X"20",X"54",X"52",
		X"49",X"47",X"47",X"45",X"52",X"20",X"20",X"20",X"52",X"49",X"47",X"48",X"54",X"20",X"54",X"52",
		X"49",X"47",X"47",X"45",X"52",X"00",X"20",X"20",X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"4D",X"41",X"43",X"48",X"49",X"4E",X"45",X"20",X"47",X"55",
		X"4E",X"20",X"00",X"20",X"4C",X"45",X"46",X"54",X"20",X"54",X"48",X"55",X"4D",X"42",X"20",X"20",
		X"20",X"20",X"20",X"52",X"49",X"47",X"48",X"54",X"20",X"54",X"48",X"55",X"4D",X"42",X"20",X"00",
		X"20",X"4F",X"49",X"4C",X"20",X"53",X"4C",X"49",X"43",X"4B",X"20",X"20",X"20",X"20",X"20",X"20",
		X"53",X"4D",X"4F",X"4B",X"45",X"20",X"53",X"43",X"52",X"45",X"45",X"4E",X"00",X"CD",X"3A",X"3D",
		X"CD",X"BC",X"89",X"21",X"5D",X"F3",X"36",X"01",X"F3",X"CD",X"93",X"01",X"FB",X"3E",X"04",X"06",
		X"90",X"21",X"70",X"E3",X"77",X"23",X"10",X"FC",X"21",X"91",X"E8",X"11",X"B5",X"96",X"CD",X"18",
		X"3F",X"21",X"DA",X"E8",X"11",X"BD",X"96",X"CD",X"18",X"3F",X"21",X"18",X"E9",X"11",X"D7",X"96",
		X"CD",X"18",X"3F",X"21",X"76",X"E9",X"11",X"ED",X"96",X"CD",X"18",X"3F",X"21",X"BA",X"E9",X"11",
		X"FF",X"96",X"CD",X"18",X"3F",X"21",X"36",X"EA",X"11",X"18",X"97",X"CD",X"18",X"3F",X"21",X"9C",
		X"EA",X"11",X"29",X"97",X"CD",X"18",X"3F",X"21",X"DC",X"EA",X"11",X"46",X"97",X"CD",X"18",X"3F",
		X"21",X"3C",X"EB",X"11",X"63",X"97",X"CD",X"18",X"3F",X"21",X"7C",X"EB",X"11",X"80",X"97",X"CD",
		X"18",X"3F",X"06",X"FF",X"CD",X"BC",X"89",X"10",X"FB",X"3E",X"FF",X"32",X"2A",X"F4",X"C9",X"03",
		X"20",X"43",X"4F",X"50",X"59",X"52",X"49",X"47",X"48",X"54",X"20",X"31",X"39",X"38",X"33",X"00",
		X"20",X"42",X"41",X"4C",X"4C",X"59",X"2F",X"4D",X"49",X"44",X"57",X"41",X"59",X"20",X"4D",X"46",
		X"47",X"20",X"43",X"4F",X"00",X"20",X"41",X"4C",X"4C",X"20",X"52",X"49",X"47",X"48",X"54",X"53",
		X"20",X"52",X"45",X"53",X"45",X"52",X"56",X"45",X"44",X"00",X"CD",X"BC",X"89",X"21",X"5D",X"F3",
		X"CD",X"2E",X"3D",X"CD",X"3A",X"3D",X"CD",X"BC",X"89",X"21",X"5D",X"F3",X"36",X"01",X"F3",X"CD",
		X"93",X"01",X"FB",X"FD",X"21",X"74",X"F8",X"FD",X"36",X"02",X"0E",X"FD",X"21",X"04",X"F8",X"11",
		X"04",X"00",X"FD",X"36",X"00",X"7C",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"1E",X"FD",X"36",
		X"03",X"68",X"FD",X"19",X"FD",X"36",X"00",X"7A",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"1F",
		X"FD",X"36",X"03",X"6D",X"FD",X"19",X"FD",X"36",X"00",X"88",X"FD",X"36",X"01",X"00",X"FD",X"36",
		X"02",X"1F",X"FD",X"36",X"03",X"68",X"FD",X"19",X"FD",X"36",X"00",X"87",X"FD",X"36",X"01",X"10",
		X"FD",X"36",X"02",X"1E",X"FD",X"36",X"03",X"6C",X"FD",X"21",X"A8",X"F8",X"FD",X"36",X"02",X"25",
		X"FD",X"36",X"06",X"00",X"3E",X"82",X"FD",X"77",X"00",X"FD",X"77",X"04",X"FD",X"36",X"03",X"F8",
		X"3E",X"E8",X"32",X"E2",X"F0",X"AF",X"FD",X"77",X"01",X"FD",X"77",X"05",X"32",X"4A",X"F0",X"32",
		X"4B",X"F0",X"32",X"4C",X"F0",X"D6",X"02",X"32",X"44",X"F0",X"CD",X"BC",X"89",X"CD",X"C9",X"9A",
		X"FD",X"7E",X"03",X"FE",X"C0",X"30",X"F3",X"3E",X"01",X"32",X"4A",X"F0",X"06",X"03",X"CD",X"BC",
		X"89",X"CD",X"C9",X"9A",X"10",X"F8",X"3E",X"01",X"32",X"4C",X"F0",X"06",X"04",X"CD",X"BC",X"89",
		X"CD",X"C9",X"9A",X"10",X"F8",X"AF",X"32",X"4C",X"F0",X"06",X"02",X"CD",X"BC",X"89",X"CD",X"C9",
		X"9A",X"10",X"F8",X"AF",X"32",X"4A",X"F0",X"D6",X"04",X"32",X"44",X"F0",X"CD",X"BC",X"89",X"CD",
		X"C9",X"9A",X"FD",X"7E",X"03",X"FE",X"78",X"30",X"F3",X"DD",X"21",X"6C",X"F8",X"3E",X"82",X"DD",
		X"77",X"00",X"DD",X"77",X"04",X"DD",X"36",X"02",X"21",X"DD",X"36",X"06",X"22",X"32",X"00",X"F0",
		X"3E",X"F8",X"32",X"01",X"F0",X"32",X"E4",X"F0",X"AF",X"32",X"D5",X"F0",X"32",X"E3",X"F0",X"3A",
		X"01",X"F0",X"D6",X"04",X"32",X"01",X"F0",X"4F",X"FE",X"E8",X"20",X"05",X"21",X"11",X"F0",X"36",
		X"01",X"FE",X"C0",X"20",X"05",X"21",X"D5",X"F0",X"36",X"20",X"DD",X"21",X"6C",X"F8",X"21",X"E4",
		X"F0",X"BE",X"20",X"15",X"FE",X"F0",X"28",X"08",X"36",X"F0",X"DD",X"36",X"02",X"00",X"18",X"09",
		X"36",X"F8",X"DD",X"36",X"06",X"00",X"C3",X"7E",X"9A",X"FE",X"34",X"C2",X"63",X"9A",X"FD",X"21",
		X"10",X"F8",X"11",X"04",X"00",X"FD",X"36",X"00",X"68",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",
		X"F0",X"FD",X"36",X"03",X"80",X"FD",X"19",X"FD",X"36",X"00",X"78",X"FD",X"36",X"01",X"00",X"FD",
		X"36",X"02",X"F1",X"FD",X"36",X"03",X"80",X"FD",X"19",X"FD",X"36",X"00",X"88",X"FD",X"36",X"01",
		X"00",X"FD",X"36",X"02",X"F2",X"FD",X"36",X"03",X"80",X"FD",X"19",X"FD",X"36",X"00",X"98",X"FD",
		X"36",X"01",X"00",X"FD",X"36",X"02",X"F3",X"FD",X"36",X"03",X"80",X"FD",X"19",X"FD",X"36",X"00",
		X"64",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"9C",X"FD",X"36",X"03",X"85",X"FD",X"19",X"FD",
		X"36",X"00",X"72",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"9D",X"FD",X"36",X"03",X"85",X"FD",
		X"19",X"FD",X"36",X"00",X"80",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"9E",X"FD",X"36",X"03",
		X"85",X"FD",X"19",X"FD",X"36",X"00",X"8E",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",X"9F",X"FD",
		X"36",X"03",X"85",X"FD",X"19",X"FD",X"36",X"00",X"9C",X"FD",X"36",X"01",X"00",X"FD",X"36",X"02",
		X"9C",X"FD",X"36",X"03",X"85",X"06",X"05",X"3E",X"02",X"21",X"43",X"F1",X"77",X"23",X"10",X"FC",
		X"32",X"E3",X"F0",X"79",X"DD",X"77",X"03",X"C6",X"10",X"DD",X"77",X"07",X"CD",X"4F",X"23",X"CD",
		X"BC",X"89",X"CD",X"C9",X"9A",X"CD",X"D1",X"9B",X"CD",X"1D",X"54",X"C3",X"6F",X"99",X"06",X"10",
		X"CD",X"BC",X"89",X"CD",X"D1",X"9B",X"10",X"F8",X"06",X"05",X"11",X"04",X"00",X"DD",X"21",X"20",
		X"F8",X"DD",X"36",X"00",X"00",X"DD",X"19",X"10",X"F8",X"21",X"36",X"EB",X"11",X"1F",X"98",X"CD",
		X"18",X"3F",X"21",X"78",X"EB",X"11",X"30",X"98",X"CD",X"18",X"3F",X"21",X"B8",X"EB",X"11",X"45",
		X"98",X"CD",X"18",X"3F",X"21",X"E3",X"F0",X"36",X"01",X"06",X"A0",X"CD",X"BC",X"89",X"CD",X"D1",
		X"9B",X"10",X"F8",X"F3",X"CD",X"93",X"01",X"FB",X"C9",X"3A",X"44",X"F0",X"B7",X"C8",X"FD",X"21",
		X"A8",X"F8",X"FD",X"86",X"03",X"FD",X"77",X"03",X"21",X"E2",X"F0",X"BE",X"20",X"23",X"FE",X"E8",
		X"20",X"08",X"36",X"F8",X"FD",X"36",X"06",X"26",X"18",X"17",X"FE",X"EC",X"28",X"08",X"36",X"EC",
		X"FD",X"36",X"02",X"00",X"18",X"0B",X"AF",X"FD",X"77",X"06",X"32",X"44",X"F0",X"32",X"11",X"F0",
		X"C9",X"DD",X"21",X"04",X"F8",X"FE",X"6C",X"20",X"43",X"11",X"04",X"00",X"DD",X"36",X"00",X"73",
		X"DD",X"36",X"01",X"20",X"DD",X"36",X"02",X"13",X"DD",X"19",X"DD",X"36",X"00",X"73",X"DD",X"36",
		X"01",X"20",X"DD",X"36",X"02",X"13",X"DD",X"36",X"03",X"6E",X"DD",X"19",X"DD",X"36",X"00",X"90",
		X"DD",X"36",X"02",X"13",X"DD",X"36",X"03",X"6C",X"DD",X"19",X"DD",X"36",X"00",X"90",X"DD",X"36",
		X"01",X"00",X"DD",X"36",X"02",X"13",X"DD",X"36",X"03",X"6E",X"18",X"4E",X"FE",X"5C",X"20",X"4A",
		X"11",X"04",X"00",X"DD",X"36",X"00",X"78",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"E8",X"DD",
		X"36",X"03",X"6A",X"DD",X"19",X"DD",X"36",X"00",X"88",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",
		X"E9",X"DD",X"36",X"03",X"6A",X"DD",X"19",X"DD",X"36",X"00",X"98",X"DD",X"36",X"02",X"E7",X"DD",
		X"36",X"03",X"6A",X"DD",X"19",X"DD",X"36",X"00",X"00",X"DD",X"21",X"41",X"F1",X"DD",X"36",X"00",
		X"03",X"DD",X"36",X"01",X"03",X"21",X"E3",X"F0",X"36",X"01",X"C6",X"10",X"FD",X"77",X"07",X"57",
		X"3A",X"4A",X"F0",X"DD",X"21",X"D8",X"F8",X"B7",X"20",X"04",X"DD",X"77",X"00",X"C9",X"DD",X"72",
		X"03",X"3A",X"4B",X"F0",X"B7",X"3E",X"0C",X"16",X"00",X"28",X"04",X"ED",X"44",X"16",X"20",X"FD",
		X"86",X"00",X"DD",X"77",X"00",X"DD",X"72",X"01",X"3A",X"4C",X"F0",X"C6",X"10",X"DD",X"77",X"02",
		X"C9",X"3A",X"E3",X"F0",X"FE",X"01",X"D8",X"C5",X"11",X"04",X"00",X"28",X"20",X"06",X"05",X"21",
		X"43",X"F1",X"DD",X"21",X"20",X"F8",X"35",X"28",X"0F",X"36",X"02",X"DD",X"7E",X"02",X"3C",X"FE",
		X"A0",X"38",X"02",X"3E",X"9C",X"DD",X"77",X"02",X"23",X"DD",X"19",X"10",X"E9",X"06",X"02",X"21",
		X"41",X"F1",X"DD",X"21",X"04",X"F8",X"35",X"20",X"10",X"36",X"03",X"DD",X"7E",X"02",X"C6",X"02",
		X"FE",X"F0",X"38",X"02",X"D6",X"08",X"DD",X"77",X"02",X"23",X"DD",X"19",X"10",X"E8",X"C1",X"C9",
		X"49",X"4E",X"54",X"52",X"4F",X"44",X"55",X"43",X"49",X"4E",X"47",X"00",X"54",X"48",X"45",X"20",
		X"45",X"4E",X"45",X"4D",X"59",X"20",X"41",X"47",X"45",X"4E",X"54",X"53",X"00",X"20",X"20",X"54",
		X"48",X"45",X"20",X"52",X"4F",X"41",X"44",X"20",X"4C",X"4F",X"52",X"44",X"20",X"00",X"20",X"42",
		X"55",X"4C",X"4C",X"45",X"54",X"20",X"50",X"52",X"4F",X"4F",X"46",X"20",X"42",X"55",X"4C",X"4C",
		X"59",X"00",X"20",X"20",X"53",X"57",X"49",X"54",X"43",X"48",X"20",X"42",X"4C",X"41",X"44",X"45",
		X"00",X"20",X"4E",X"45",X"56",X"45",X"52",X"20",X"54",X"4F",X"20",X"42",X"45",X"20",X"54",X"52",
		X"55",X"53",X"54",X"45",X"44",X"00",X"20",X"20",X"54",X"48",X"45",X"20",X"45",X"4E",X"46",X"4F",
		X"52",X"43",X"45",X"52",X"00",X"44",X"4F",X"55",X"42",X"4C",X"45",X"20",X"42",X"41",X"52",X"52",
		X"45",X"4C",X"20",X"41",X"43",X"54",X"49",X"4F",X"4E",X"00",X"20",X"54",X"48",X"45",X"20",X"4D",
		X"41",X"44",X"20",X"42",X"4F",X"4D",X"42",X"45",X"52",X"00",X"20",X"20",X"4D",X"41",X"53",X"54",
		X"45",X"52",X"20",X"4F",X"46",X"20",X"54",X"48",X"45",X"20",X"53",X"4B",X"59",X"00",X"41",X"56",
		X"4F",X"49",X"44",X"20",X"41",X"4C",X"4C",X"20",X"4F",X"54",X"48",X"45",X"52",X"20",X"43",X"41",
		X"52",X"53",X"00",X"20",X"20",X"41",X"4E",X"44",X"20",X"4D",X"4F",X"54",X"4F",X"52",X"43",X"59",
		X"43",X"4C",X"45",X"53",X"20",X"20",X"20",X"00",X"20",X"20",X"20",X"57",X"52",X"45",X"43",X"4B",
		X"49",X"4E",X"47",X"20",X"54",X"48",X"45",X"4D",X"20",X"20",X"20",X"20",X"00",X"54",X"45",X"4D",
		X"50",X"4F",X"52",X"41",X"52",X"49",X"4C",X"59",X"20",X"44",X"49",X"53",X"41",X"42",X"4C",X"45",
		X"53",X"00",X"20",X"20",X"20",X"50",X"4F",X"49",X"4E",X"54",X"20",X"53",X"43",X"4F",X"52",X"49",
		X"4E",X"47",X"00",X"31",X"35",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"35",X"30",
		X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"37",X"30",X"30",X"20",X"50",X"4F",X"49",
		X"4E",X"54",X"53",X"00",X"CD",X"BC",X"89",X"21",X"5D",X"F3",X"CD",X"2E",X"3D",X"CD",X"3A",X"3D",
		X"CD",X"BC",X"89",X"21",X"5D",X"F3",X"36",X"01",X"F3",X"CD",X"93",X"01",X"FB",X"AF",X"32",X"01",
		X"F4",X"CD",X"BE",X"11",X"CD",X"BC",X"89",X"AF",X"32",X"33",X"F0",X"32",X"35",X"F0",X"32",X"81",
		X"F0",X"32",X"82",X"F0",X"32",X"6C",X"F3",X"32",X"06",X"F0",X"32",X"03",X"F0",X"32",X"A1",X"F0",
		X"3C",X"32",X"01",X"F4",X"21",X"FA",X"B9",X"22",X"3C",X"F0",X"21",X"00",X"F0",X"36",X"CC",X"21",
		X"02",X"F0",X"36",X"08",X"21",X"93",X"E8",X"11",X"20",X"9C",X"CD",X"18",X"3F",X"21",X"D6",X"E8",
		X"11",X"2C",X"9C",X"CD",X"18",X"3F",X"CD",X"BC",X"89",X"CD",X"DF",X"8B",X"3A",X"03",X"F0",X"B7",
		X"20",X"39",X"3A",X"00",X"F0",X"D6",X"84",X"28",X"06",X"3E",X"01",X"30",X"02",X"ED",X"44",X"32",
		X"A1",X"F0",X"AF",X"32",X"06",X"F0",X"3A",X"82",X"F0",X"FE",X"0A",X"06",X"20",X"3A",X"81",X"F0",
		X"20",X"05",X"B7",X"28",X"16",X"06",X"01",X"21",X"82",X"F0",X"38",X"06",X"90",X"30",X"07",X"35",
		X"18",X"04",X"80",X"30",X"01",X"34",X"32",X"81",X"F0",X"18",X"BB",X"3A",X"6C",X"F3",X"47",X"CB",
		X"27",X"80",X"21",X"0B",X"9E",X"85",X"30",X"01",X"24",X"6F",X"E9",X"C3",X"32",X"9E",X"C3",X"68",
		X"9E",X"C3",X"84",X"9E",X"C3",X"68",X"9E",X"C3",X"B9",X"9E",X"C3",X"F4",X"9E",X"C3",X"FE",X"9E",
		X"C3",X"68",X"9E",X"C3",X"16",X"9F",X"C3",X"68",X"9E",X"C3",X"46",X"9F",X"C3",X"51",X"9F",X"C3",
		X"E8",X"9F",X"DD",X"21",X"8B",X"F2",X"DD",X"7E",X"01",X"B7",X"C2",X"B6",X"9D",X"CD",X"58",X"0D",
		X"21",X"93",X"E8",X"CD",X"15",X"3F",X"21",X"D6",X"E8",X"11",X"3D",X"9C",X"CD",X"18",X"3F",X"21",
		X"58",X"EB",X"11",X"4E",X"9C",X"CD",X"18",X"3F",X"21",X"93",X"EB",X"11",X"33",X"9D",X"CD",X"18",
		X"3F",X"21",X"6C",X"F3",X"34",X"C3",X"B6",X"9D",X"3A",X"03",X"F0",X"E6",X"01",X"CA",X"B6",X"9D",
		X"21",X"D6",X"E8",X"CD",X"15",X"3F",X"21",X"58",X"EB",X"CD",X"15",X"3F",X"21",X"98",X"EB",X"CD",
		X"15",X"3F",X"18",X"DD",X"3A",X"82",X"F0",X"FE",X"0A",X"C2",X"B6",X"9D",X"DD",X"21",X"8B",X"F2",
		X"DD",X"7E",X"01",X"B7",X"C2",X"B6",X"9D",X"3E",X"03",X"CD",X"58",X"0D",X"21",X"D6",X"E8",X"11",
		X"62",X"9C",X"CD",X"18",X"3F",X"21",X"58",X"EB",X"11",X"71",X"9C",X"CD",X"18",X"3F",X"21",X"93",
		X"EB",X"11",X"33",X"9D",X"CD",X"18",X"3F",X"18",X"A8",X"3A",X"82",X"F0",X"FE",X"0A",X"C2",X"B6",
		X"9D",X"DD",X"21",X"8B",X"F2",X"DD",X"7E",X"01",X"B7",X"C2",X"B6",X"9D",X"3C",X"32",X"45",X"F0",
		X"32",X"42",X"F0",X"CD",X"76",X"0C",X"21",X"D6",X"E8",X"11",X"86",X"9C",X"CD",X"18",X"3F",X"21",
		X"58",X"EB",X"11",X"95",X"9C",X"CD",X"18",X"3F",X"21",X"93",X"EB",X"11",X"3E",X"9D",X"CD",X"18",
		X"3F",X"C3",X"61",X"9E",X"3A",X"42",X"F0",X"B7",X"C2",X"B6",X"9D",X"C3",X"61",X"9E",X"DD",X"21",
		X"8B",X"F2",X"DD",X"7E",X"01",X"B7",X"C2",X"B6",X"9D",X"32",X"2F",X"F0",X"3C",X"32",X"45",X"F0",
		X"CD",X"76",X"0C",X"C3",X"61",X"9E",X"3A",X"00",X"F0",X"FE",X"84",X"C2",X"B6",X"9D",X"21",X"FC",
		X"F0",X"36",X"0A",X"21",X"E8",X"F0",X"36",X"01",X"21",X"D6",X"E8",X"11",X"AA",X"9C",X"CD",X"18",
		X"3F",X"21",X"58",X"EB",X"11",X"BA",X"9C",X"CD",X"18",X"3F",X"21",X"93",X"EB",X"11",X"49",X"9D",
		X"CD",X"18",X"3F",X"C3",X"61",X"9E",X"3A",X"82",X"F0",X"FE",X"0A",X"C2",X"B6",X"9D",X"C3",X"61",
		X"9E",X"DD",X"21",X"8B",X"F2",X"11",X"23",X"00",X"06",X"06",X"DD",X"7E",X"01",X"B7",X"28",X"07",
		X"DD",X"19",X"10",X"F6",X"C3",X"B6",X"9D",X"DD",X"22",X"48",X"F0",X"21",X"D9",X"B9",X"22",X"3C",
		X"F0",X"3A",X"00",X"F0",X"DD",X"77",X"05",X"3A",X"01",X"F0",X"DD",X"77",X"07",X"DD",X"36",X"02",
		X"14",X"DD",X"36",X"06",X"21",X"DD",X"36",X"1D",X"22",X"DD",X"36",X"0E",X"14",X"DD",X"36",X"0F",
		X"03",X"DD",X"36",X"03",X"0A",X"DD",X"36",X"0B",X"0C",X"DD",X"36",X"01",X"80",X"DD",X"36",X"0C",
		X"01",X"AF",X"DD",X"77",X"08",X"DD",X"77",X"1F",X"DD",X"77",X"0A",X"DD",X"77",X"10",X"DD",X"77",
		X"04",X"32",X"00",X"F0",X"32",X"01",X"F0",X"3E",X"04",X"32",X"33",X"F0",X"32",X"35",X"F0",X"21",
		X"03",X"F0",X"36",X"90",X"21",X"06",X"F0",X"36",X"02",X"21",X"6D",X"F3",X"36",X"FF",X"21",X"2F",
		X"F0",X"36",X"03",X"21",X"98",X"E8",X"11",X"CE",X"9C",X"CD",X"18",X"3F",X"21",X"D8",X"E8",X"11",
		X"E3",X"9C",X"CD",X"18",X"3F",X"C3",X"61",X"9E",X"DD",X"2A",X"48",X"F0",X"21",X"82",X"F0",X"DD",
		X"4E",X"03",X"DD",X"7E",X"07",X"FE",X"68",X"38",X"07",X"FE",X"D0",X"38",X"05",X"0D",X"18",X"02",
		X"00",X"00",X"00",X"0F",X"CC",X"03",X"00",X"2B",X"C4",X"0F",X"01",X"00",X"00",X"77",X"CC",X"04",
		X"00",X"67",X"C4",X"0F",X"00",X"00",X"00",X"D7",X"CC",X"04",X"00",X"67",X"C4",X"03",X"00",X"6B",
		X"C4",X"0B",X"00",X"00",X"00",X"23",X"CD",X"04",X"00",X"6B",X"C4",X"0F",X"00",X"00",X"00",X"63",
		X"CD",X"04",X"00",X"6B",X"C4",X"0B",X"00",X"67",X"C4",X"03",X"00",X"00",X"00",X"AF",X"CD",X"03",
		X"00",X"6F",X"C4",X"0E",X"01",X"27",X"C4",X"00",X"00",X"17",X"CE",X"03",X"00",X"AB",X"C4",X"0F",
		X"01",X"00",X"00",X"7F",X"CE",X"04",X"00",X"E7",X"C4",X"0F",X"00",X"00",X"00",X"DF",X"CE",X"04",
		X"00",X"E7",X"C4",X"03",X"00",X"EB",X"C4",X"0B",X"00",X"00",X"00",X"2B",X"CF",X"04",X"00",X"EB",
		X"C4",X"0F",X"00",X"00",X"00",X"6B",X"CF",X"04",X"00",X"EB",X"C4",X"0B",X"00",X"E7",X"C4",X"03",
		X"00",X"00",X"00",X"E4",X"CF",X"03",X"00",X"EF",X"C4",X"0E",X"01",X"27",X"C4",X"00",X"00",X"4C",
		X"D0",X"04",X"00",X"27",X"C4",X"03",X"00",X"2B",X"C5",X"0B",X"00",X"00",X"00",X"A2",X"D0",X"04",
		X"00",X"2B",X"C5",X"0F",X"00",X"00",X"00",X"F2",X"D0",X"04",X"00",X"2B",X"C5",X"0B",X"00",X"27",
		X"C4",X"03",X"00",X"00",X"00",X"48",X"D1",X"05",X"00",X"27",X"C4",X"17",X"C4",X"13",X"C4",X"0B",
		X"C4",X"03",X"C4",X"FB",X"C3",X"F7",X"C3",X"F3",X"C3",X"EF",X"C3",X"EB",X"C3",X"DF",X"C3",X"D7",
		X"C3",X"CB",X"C3",X"C7",X"C3",X"BF",X"C3",X"BB",X"C3",X"00",X"00",X"A0",X"D1",X"05",X"00",X"2F",
		X"C5",X"0F",X"01",X"00",X"00",X"EC",X"D1",X"05",X"00",X"6F",X"C5",X"0F",X"00",X"00",X"00",X"34",
		X"D2",X"04",X"00",X"6F",X"C5",X"0F",X"01",X"00",X"00",X"8A",X"D2",X"04",X"00",X"AF",X"C5",X"03",
		X"00",X"B3",X"C5",X"0B",X"00",X"00",X"00",X"E2",X"D2",X"04",X"00",X"B3",X"C5",X"0F",X"00",X"00",
		X"00",X"3A",X"D3",X"04",X"00",X"AF",X"C5",X"03",X"00",X"A3",X"C5",X"9B",X"C5",X"93",X"C5",X"8B",
		X"C5",X"83",X"C5",X"7B",X"C5",X"77",X"C5",X"73",X"C5",X"6F",X"C5",X"03",X"00",X"00",X"00",X"8E",
		X"D3",X"04",X"00",X"6F",X"C5",X"04",X"00",X"B7",X"C5",X"0A",X"01",X"00",X"00",X"E0",X"D3",X"05",
		X"00",X"DF",X"C5",X"DF",X"C5",X"0E",X"01",X"00",X"00",X"3A",X"D4",X"05",X"00",X"1B",X"C6",X"0D",
		X"01",X"B3",X"C3",X"B3",X"C3",X"00",X"00",X"83",X"D4",X"05",X"00",X"DF",X"C5",X"DF",X"C5",X"53",
		X"C6",X"0D",X"01",X"00",X"00",X"DD",X"D4",X"05",X"00",X"8B",X"C6",X"0C",X"01",X"B3",X"C3",X"02",
		X"00",X"00",X"00",X"26",X"D5",X"04",X"00",X"E7",X"C4",X"BF",X"C6",X"0E",X"01",X"00",X"00",X"7E",
		X"D5",X"04",X"00",X"FB",X"C6",X"0F",X"01",X"00",X"00",X"D5",X"D5",X"01",X"00",X"3B",X"C7",X"3B",
		X"C7",X"3F",X"C7",X"3F",X"C7",X"43",X"C7",X"43",X"C7",X"47",X"C7",X"47",X"C7",X"4B",X"C7",X"03",
		X"01",X"5B",X"C7",X"5B",X"C7",X"5F",X"C7",X"63",X"C7",X"00",X"00",X"35",X"D6",X"01",X"00",X"67",
		X"C7",X"02",X"01",X"73",X"C7",X"02",X"00",X"77",X"C7",X"03",X"00",X"EB",X"C4",X"05",X"00",X"00",
		X"00",X"7D",X"D6",X"04",X"00",X"EB",X"C4",X"0B",X"00",X"E7",X"C4",X"03",X"00",X"00",X"00",X"C5",
		X"D6",X"04",X"00",X"E7",X"C4",X"0F",X"00",X"00",X"00",X"23",X"D7",X"04",X"00",X"E7",X"C4",X"0F",
		X"00",X"00",X"00",X"C6",X"D7",X"01",X"00",X"7F",X"C7",X"0F",X"00",X"00",X"00",X"F6",X"D7",X"01",
		X"00",X"8F",X"C7",X"07",X"00",X"93",X"C7",X"97",X"C7",X"9B",X"C7",X"05",X"00",X"00",X"00",X"3B",
		X"D8",X"01",X"00",X"9B",X"C7",X"03",X"00",X"9F",X"C7",X"0B",X"00",X"00",X"00",X"91",X"D8",X"01",
		X"00",X"9F",X"C7",X"0F",X"00",X"00",X"00",X"E9",X"D8",X"01",X"00",X"9F",X"C7",X"05",X"00",X"A3",
		X"C7",X"05",X"00",X"9B",X"C7",X"03",X"00",X"00",X"00",X"4B",X"D9",X"01",X"00",X"9B",X"C7",X"03",
		X"00",X"A7",X"C7",X"9F",X"C7",X"06",X"00",X"9B",X"C7",X"03",X"00",X"00",X"00",X"9F",X"D9",X"01",
		X"00",X"63",X"C8",X"63",X"C8",X"AB",X"C7",X"04",X"01",X"BB",X"C7",X"03",X"01",X"9F",X"C7",X"04",
		X"00",X"00",X"00",X"05",X"DA",X"01",X"00",X"9F",X"C7",X"9F",X"C7",X"CB",X"C7",X"CF",X"C7",X"02",
		X"00",X"D3",X"C7",X"02",X"01",X"8F",X"C7",X"02",X"01",X"9B",X"C7",X"03",X"00",X"00",X"00",X"09",
		X"DE",X"01",X"00",X"63",X"C8",X"04",X"00",X"FF",X"C7",X"0A",X"01",X"00",X"00",X"58",X"DA",X"01",
		X"00",X"FF",X"C8",X"FF",X"C8",X"DF",X"C7",X"DF",X"C7",X"E3",X"C7",X"E3",X"C7",X"F7",X"C7",X"04",
		X"00",X"E7",X"C7",X"04",X"00",X"00",X"00",X"BB",X"DA",X"01",X"00",X"E7",X"C7",X"E7",X"C7",X"EB",
		X"C7",X"EB",X"C7",X"EF",X"C7",X"EB",X"C7",X"EB",X"C7",X"F3",X"C7",X"08",X"00",X"00",X"00",X"24",
		X"DB",X"01",X"00",X"F3",X"C7",X"08",X"00",X"4B",X"C8",X"06",X"00",X"00",X"00",X"8C",X"DB",X"01",
		X"00",X"4B",X"C8",X"4B",X"C8",X"4F",X"C8",X"03",X"00",X"53",X"C8",X"09",X"00",X"00",X"00",X"E8",
		X"DB",X"02",X"00",X"57",X"C8",X"0F",X"00",X"00",X"00",X"38",X"DC",X"02",X"00",X"57",X"C8",X"03",
		X"00",X"5B",X"C8",X"5F",X"C8",X"5F",X"C8",X"5B",X"C8",X"63",X"C8",X"63",X"C8",X"67",X"C8",X"02",
		X"00",X"63",X"C8",X"02",X"00",X"00",X"00",X"94",X"DC",X"02",X"00",X"63",X"C8",X"0F",X"00",X"00",
		X"00",X"DC",X"DC",X"02",X"00",X"63",X"C8",X"04",X"00",X"6B",X"C8",X"6F",X"C8",X"09",X"00",X"00",
		X"00",X"1F",X"DD",X"02",X"00",X"6F",X"C8",X"0F",X"00",X"00",X"00",X"5F",X"DD",X"01",X"00",X"9B",
		X"C7",X"05",X"00",X"63",X"C8",X"09",X"00",X"00",X"00",X"AA",X"DD",X"01",X"00",X"6F",X"C8",X"73",
		X"C8",X"77",X"C8",X"77",X"C8",X"7B",X"C8",X"03",X"00",X"9B",X"C7",X"03",X"00",X"7F",X"C8",X"83",
		X"C8",X"02",X"00",X"00",X"00",X"7D",X"DE",X"01",X"00",X"E7",X"C4",X"0F",X"00",X"00",X"00",X"DD",
		X"DE",X"03",X"00",X"2B",X"C8",X"02",X"00",X"6F",X"C7",X"2F",X"C8",X"2F",X"C8",X"33",X"C8",X"33",
		X"C8",X"37",X"C8",X"3B",X"C8",X"3F",X"C8",X"3F",X"C8",X"43",X"C8",X"47",X"C8",X"87",X"C8",X"8B",
		X"C8",X"00",X"00",X"3D",X"DF",X"04",X"00",X"8F",X"C8",X"0F",X"01",X"00",X"00",X"98",X"DF",X"04",
		X"00",X"CF",X"C8",X"E7",X"C4",X"0E",X"00",X"00",X"00",X"45",X"DE",X"01",X"00",X"D3",X"C8",X"0A",
		X"01",X"FF",X"C8",X"04",X"00",X"00",X"00",X"83",X"D7",X"01",X"00",X"7F",X"C7",X"0F",X"00",X"00",
		X"00",X"B7",X"CF",X"04",X"00",X"EB",X"C4",X"03",X"00",X"7B",X"C7",X"07",X"00",X"EB",X"C4",X"03",
		X"00",X"00",X"00",X"02",X"32",X"92",X"00",X"02",X"33",X"91",X"00",X"02",X"34",X"8F",X"00",X"02",
		X"35",X"8D",X"00",X"02",X"36",X"8B",X"00",X"02",X"37",X"88",X"00",X"02",X"38",X"84",X"00",X"02",
		X"39",X"82",X"00",X"02",X"3A",X"80",X"00",X"02",X"3B",X"7F",X"00",X"02",X"3D",X"7D",X"00",X"02",
		X"3D",X"7C",X"00",X"02",X"3E",X"7A",X"00",X"02",X"40",X"78",X"00",X"02",X"40",X"75",X"00",X"02",
		X"42",X"72",X"00",X"02",X"43",X"70",X"00",X"02",X"45",X"6C",X"00",X"02",X"47",X"68",X"00",X"02",
		X"47",X"67",X"00",X"02",X"49",X"65",X"00",X"02",X"4A",X"64",X"00",X"02",X"4B",X"60",X"00",X"02",
		X"4C",X"5E",X"00",X"02",X"4D",X"5C",X"00",X"02",X"50",X"56",X"00",X"02",X"50",X"54",X"00",X"02",
		X"51",X"52",X"00",X"02",X"52",X"51",X"00",X"02",X"52",X"50",X"00",X"42",X"50",X"50",X"00",X"42",
		X"4C",X"52",X"00",X"42",X"4B",X"53",X"00",X"42",X"49",X"52",X"00",X"42",X"45",X"52",X"00",X"42",
		X"41",X"52",X"00",X"42",X"3C",X"52",X"00",X"42",X"38",X"52",X"00",X"42",X"34",X"52",X"00",X"42",
		X"32",X"51",X"00",X"42",X"30",X"4D",X"00",X"42",X"2C",X"4D",X"00",X"42",X"2B",X"4C",X"00",X"42",
		X"29",X"4B",X"00",X"42",X"26",X"4D",X"00",X"02",X"24",X"4F",X"00",X"82",X"24",X"4F",X"00",X"22",
		X"23",X"52",X"00",X"22",X"24",X"52",X"00",X"22",X"27",X"52",X"00",X"22",X"2A",X"52",X"00",X"22",
		X"2D",X"52",X"00",X"22",X"31",X"52",X"00",X"22",X"35",X"52",X"00",X"22",X"39",X"53",X"00",X"22",
		X"3D",X"54",X"00",X"22",X"41",X"53",X"00",X"22",X"46",X"51",X"00",X"22",X"4A",X"4F",X"00",X"22",
		X"4E",X"4D",X"00",X"22",X"51",X"4D",X"00",X"22",X"52",X"4E",X"00",X"22",X"52",X"54",X"00",X"22",
		X"53",X"54",X"00",X"22",X"55",X"55",X"00",X"22",X"57",X"55",X"00",X"22",X"5D",X"53",X"00",X"22",
		X"61",X"55",X"00",X"22",X"65",X"55",X"00",X"22",X"68",X"58",X"00",X"22",X"6C",X"57",X"00",X"22",
		X"71",X"54",X"00",X"22",X"75",X"52",X"00",X"22",X"7A",X"50",X"00",X"22",X"7E",X"4D",X"00",X"22",
		X"81",X"4C",X"00",X"22",X"82",X"4D",X"00",X"02",X"82",X"50",X"00",X"82",X"82",X"50",X"00",X"42",
		X"80",X"52",X"00",X"42",X"7C",X"52",X"00",X"42",X"7A",X"54",X"00",X"42",X"78",X"54",X"00",X"42",
		X"75",X"53",X"00",X"42",X"6F",X"54",X"00",X"42",X"6B",X"55",X"00",X"42",X"66",X"56",X"00",X"42",
		X"63",X"55",X"00",X"42",X"60",X"53",X"00",X"42",X"5E",X"52",X"00",X"42",X"5C",X"50",X"00",X"42",
		X"5A",X"4E",X"00",X"42",X"58",X"4C",X"00",X"42",X"55",X"4E",X"00",X"82",X"52",X"50",X"00",X"02",
		X"31",X"93",X"00",X"02",X"2F",X"97",X"00",X"02",X"2D",X"9B",X"00",X"02",X"2B",X"9F",X"00",X"02",
		X"28",X"A4",X"00",X"02",X"26",X"A8",X"00",X"02",X"24",X"AC",X"00",X"04",X"22",X"B0",X"00",X"04",
		X"22",X"50",X"12",X"04",X"20",X"50",X"16",X"04",X"1D",X"4F",X"1B",X"04",X"1B",X"4F",X"20",X"04",
		X"19",X"50",X"22",X"04",X"17",X"50",X"25",X"04",X"15",X"52",X"27",X"04",X"14",X"51",X"2B",X"05",
		X"12",X"50",X"10",X"05",X"12",X"4F",X"14",X"05",X"12",X"4D",X"18",X"05",X"12",X"4C",X"1A",X"05",
		X"12",X"4B",X"1C",X"05",X"12",X"4A",X"1E",X"05",X"12",X"49",X"20",X"05",X"12",X"48",X"22",X"05",
		X"12",X"47",X"24",X"05",X"12",X"46",X"26",X"05",X"12",X"45",X"28",X"05",X"12",X"44",X"2A",X"05",
		X"12",X"43",X"2C",X"05",X"12",X"42",X"2E",X"05",X"12",X"41",X"30",X"05",X"12",X"40",X"32",X"05",
		X"12",X"40",X"31",X"85",X"12",X"40",X"30",X"05",X"14",X"4E",X"10",X"05",X"15",X"4D",X"10",X"05",
		X"17",X"4B",X"10",X"05",X"18",X"4A",X"10",X"05",X"19",X"49",X"10",X"05",X"1A",X"4C",X"0A",X"05",
		X"1B",X"4D",X"06",X"05",X"1C",X"4E",X"02",X"05",X"1D",X"4D",X"02",X"05",X"1F",X"4B",X"02",X"05",
		X"21",X"49",X"02",X"05",X"26",X"48",X"05",X"05",X"2B",X"47",X"04",X"05",X"2F",X"47",X"04",X"05",
		X"31",X"47",X"04",X"05",X"32",X"47",X"06",X"05",X"32",X"49",X"05",X"07",X"32",X"4B",X"07",X"07",
		X"32",X"4F",X"08",X"07",X"32",X"52",X"08",X"07",X"32",X"56",X"07",X"07",X"32",X"5A",X"08",X"07",
		X"32",X"5E",X"07",X"07",X"32",X"62",X"07",X"07",X"32",X"66",X"08",X"07",X"32",X"6A",X"08",X"07",
		X"32",X"6E",X"08",X"07",X"32",X"72",X"08",X"07",X"32",X"76",X"08",X"07",X"32",X"7A",X"08",X"07",
		X"32",X"7E",X"08",X"07",X"32",X"82",X"08",X"07",X"32",X"86",X"08",X"07",X"32",X"8A",X"08",X"07",
		X"32",X"8E",X"08",X"07",X"32",X"92",X"08",X"07",X"32",X"92",X"09",X"07",X"32",X"92",X"0A",X"07",
		X"32",X"92",X"0B",X"05",X"1C",X"48",X"05",X"05",X"19",X"47",X"04",X"05",X"15",X"47",X"04",X"05",
		X"13",X"47",X"04",X"05",X"10",X"47",X"06",X"05",X"0B",X"49",X"05",X"06",X"52",X"07",X"4B",X"06",
		X"4E",X"08",X"4E",X"06",X"4A",X"08",X"52",X"06",X"46",X"07",X"57",X"06",X"42",X"08",X"5A",X"06",
		X"3E",X"07",X"60",X"06",X"3A",X"07",X"63",X"06",X"36",X"08",X"66",X"06",X"32",X"08",X"6A",X"06",
		X"2E",X"08",X"6E",X"06",X"2A",X"08",X"72",X"06",X"22",X"08",X"76",X"06",X"1E",X"08",X"7A",X"06",
		X"1A",X"08",X"7E",X"06",X"16",X"08",X"82",X"06",X"12",X"08",X"86",X"06",X"0E",X"08",X"8A",X"06",
		X"0A",X"08",X"8E",X"06",X"06",X"08",X"92",X"06",X"02",X"0C",X"92",X"06",X"01",X"0D",X"92",X"01",
		X"80",X"02",X"50",X"01",X"7E",X"04",X"50",X"01",X"7C",X"06",X"50",X"01",X"7A",X"08",X"50",X"01",
		X"77",X"0B",X"50",X"01",X"73",X"0F",X"50",X"01",X"6D",X"15",X"50",X"01",X"68",X"1A",X"50",X"01",
		X"64",X"1E",X"50",X"01",X"62",X"20",X"50",X"01",X"60",X"22",X"50",X"01",X"5E",X"24",X"50",X"01",
		X"5C",X"26",X"50",X"01",X"5A",X"28",X"50",X"01",X"56",X"2C",X"50",X"01",X"53",X"2F",X"50",X"01",
		X"50",X"32",X"50",X"01",X"4E",X"34",X"50",X"01",X"4C",X"36",X"50",X"01",X"48",X"3A",X"50",X"01",
		X"44",X"3E",X"50",X"08",X"40",X"24",X"60",X"08",X"3B",X"29",X"60",X"08",X"36",X"2E",X"60",X"09",
		X"32",X"2A",X"58",X"09",X"2F",X"2B",X"58",X"03",X"2D",X"2F",X"08",X"03",X"2B",X"29",X"10",X"03",
		X"2A",X"26",X"14",X"03",X"28",X"24",X"18",X"03",X"26",X"23",X"1B",X"03",X"24",X"22",X"1E",X"03",
		X"24",X"20",X"20",X"03",X"24",X"1F",X"21",X"03",X"24",X"1E",X"22",X"03",X"24",X"1C",X"24",X"03",
		X"24",X"1A",X"26",X"0F",X"24",X"18",X"28",X"03",X"24",X"16",X"2A",X"03",X"24",X"15",X"2B",X"03",
		X"24",X"14",X"2C",X"03",X"24",X"13",X"2D",X"03",X"24",X"12",X"2E",X"03",X"24",X"11",X"2F",X"03",
		X"24",X"10",X"30",X"03",X"21",X"14",X"2F",X"00",X"29",X"04",X"37",X"8E",X"00",X"00",X"00",X"02",
		X"40",X"A8",X"00",X"02",X"38",X"A8",X"00",X"02",X"3C",X"A4",X"00",X"02",X"40",X"A0",X"00",X"02",
		X"44",X"90",X"00",X"02",X"44",X"88",X"00",X"02",X"44",X"80",X"00",X"02",X"44",X"70",X"00",X"02",
		X"44",X"60",X"00",X"04",X"44",X"20",X"20",X"02",X"44",X"68",X"00",X"0B",X"24",X"3C",X"50",X"0C",
		X"2C",X"38",X"38",X"0D",X"18",X"28",X"28",X"0D",X"18",X"28",X"28",X"0D",X"20",X"20",X"20",X"0C",
		X"20",X"38",X"28",X"0B",X"20",X"40",X"30",X"02",X"30",X"70",X"00",X"02",X"44",X"50",X"00",X"02",
		X"44",X"40",X"00",X"0D",X"44",X"40",X"1C",X"0C",X"44",X"50",X"28",X"02",X"44",X"98",X"00",X"09",
		X"22",X"3E",X"44",X"0A",X"22",X"32",X"30",X"0A",X"32",X"2C",X"26",X"0A",X"32",X"32",X"1C",X"00",
		X"32",X"32",X"1C",X"02",X"32",X"42",X"00",X"0F",X"26",X"28",X"2C",X"0F",X"2C",X"32",X"26",X"01",
		X"24",X"90",X"08",X"01",X"24",X"90",X"10",X"01",X"24",X"8C",X"14",X"01",X"24",X"88",X"18",X"01",
		X"24",X"84",X"1C",X"01",X"24",X"80",X"20",X"01",X"24",X"7C",X"24",X"01",X"24",X"78",X"28",X"01",
		X"24",X"74",X"2C",X"01",X"24",X"70",X"30",X"01",X"24",X"6C",X"34",X"03",X"22",X"12",X"30",X"03",
		X"26",X"12",X"26",X"03",X"28",X"12",X"2A",X"03",X"28",X"16",X"26",X"03",X"2A",X"16",X"24",X"03",
		X"2C",X"18",X"20",X"03",X"2E",X"18",X"1E",X"03",X"32",X"10",X"1A",X"02",X"34",X"40",X"00",X"02",
		X"34",X"50",X"00",X"02",X"34",X"60",X"00",X"02",X"34",X"70",X"00",X"0B",X"34",X"28",X"38",X"0C",
		X"34",X"20",X"30",X"02",X"34",X"80",X"00",X"0C",X"34",X"40",X"28",X"02",X"34",X"88",X"00",X"02",
		X"34",X"90",X"00",X"0B",X"34",X"38",X"48",X"0C",X"34",X"30",X"40",X"0C",X"44",X"20",X"40",X"0B",
		X"44",X"38",X"28",X"0C",X"44",X"30",X"20",X"03",X"36",X"18",X"16",X"03",X"3A",X"18",X"12",X"03",
		X"3E",X"18",X"0E",X"03",X"42",X"18",X"0A",X"03",X"46",X"18",X"06",X"03",X"4A",X"18",X"02",X"08",
		X"4E",X"16",X"50",X"09",X"52",X"18",X"58",X"01",X"56",X"24",X"58",X"01",X"5A",X"20",X"58",X"01",
		X"5E",X"1C",X"58",X"01",X"62",X"18",X"58",X"01",X"66",X"12",X"58",X"01",X"6A",X"0E",X"58",X"01",
		X"6E",X"0A",X"58",X"01",X"72",X"06",X"58",X"01",X"76",X"02",X"58",X"02",X"7A",X"58",X"00",X"02",
		X"7E",X"54",X"00",X"01",X"24",X"68",X"38",X"01",X"24",X"64",X"3C",X"01",X"24",X"60",X"40",X"01",
		X"24",X"5C",X"44",X"01",X"24",X"58",X"48",X"01",X"24",X"54",X"4C",X"01",X"24",X"50",X"50",X"01",
		X"24",X"4C",X"54",X"01",X"24",X"4A",X"56",X"01",X"24",X"48",X"58",X"01",X"24",X"46",X"5A",X"01",
		X"24",X"44",X"5C",X"00",X"DB",X"01",X"81",X"01",X"01",X"00",X"92",X"01",X"D0",X"01",X"6D",X"01",
		X"C7",X"01",X"E8",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"7C",X"00",X"03",X"01",X"30",X"00",
		X"1B",X"01",X"FF",X"00",X"49",X"01",X"CE",X"00",X"A9",X"00",X"07",X"01",X"80",X"01",X"4B",X"00",
		X"2B",X"00",X"04",X"01",X"52",X"00",X"00",X"00",X"21",X"00",X"02",X"01",X"24",X"00",X"13",X"01",
		X"01",X"01",X"FF",X"00",X"49",X"01",X"CE",X"00",X"A9",X"01",X"C6",X"01",X"80",X"01",X"1C",X"00",
		X"2B",X"01",X"4B",X"01",X"52",X"00",X"00",X"00",X"21",X"01",X"01",X"01",X"24",X"00",X"13",X"01",
		X"01",X"01",X"FF",X"00",X"49",X"01",X"CE",X"00",X"A9",X"01",X"5F",X"01",X"80",X"01",X"13",X"00",
		X"2B",X"01",X"1C",X"01",X"52",X"00",X"00",X"00",X"21",X"00",X"02",X"01",X"24",X"00",X"13",X"01",
		X"01",X"01",X"FF",X"01",X"24",X"01",X"CE",X"00",X"A9",X"00",X"34",X"01",X"80",X"00",X"DB",X"00",
		X"2B",X"01",X"6D",X"01",X"52",X"00",X"00",X"00",X"21",X"00",X"22",X"01",X"24",X"00",X"13",X"00",
		X"92",X"01",X"FF",X"00",X"49",X"01",X"CE",X"00",X"A9",X"00",X"90",X"01",X"80",X"01",X"1C",X"00",
		X"2B",X"01",X"13",X"01",X"52",X"00",X"00",X"00",X"21",X"01",X"01",X"01",X"24",X"00",X"13",X"00",
		X"92",X"01",X"FF",X"00",X"49",X"01",X"CE",X"00",X"A9",X"01",X"1E",X"01",X"80",X"01",X"13",X"00",
		X"2B",X"00",X"14",X"01",X"52",X"00",X"00",X"00",X"21",X"00",X"02",X"01",X"24",X"00",X"13",X"01",
		X"01",X"01",X"FF",X"02",X"40",X"C1",X"44",X"09",X"81",X"00",X"02",X"02",X"41",X"C1",X"44",X"09",
		X"81",X"41",X"02",X"42",X"00",X"C1",X"44",X"09",X"81",X"01",X"02",X"02",X"01",X"C1",X"44",X"09",
		X"81",X"40",X"02",X"02",X"40",X"C1",X"44",X"09",X"81",X"41",X"02",X"02",X"41",X"C1",X"44",X"09",
		X"81",X"00",X"02",X"02",X"00",X"C1",X"44",X"09",X"81",X"01",X"02",X"02",X"01",X"C1",X"44",X"09",
		X"81",X"40",X"02",X"02",X"41",X"C1",X"44",X"09",X"81",X"40",X"02",X"02",X"40",X"C1",X"44",X"09",
		X"81",X"02",X"41",X"AD",X"02",X"C1",X"44",X"09",X"81",X"01",X"02",X"02",X"41",X"C1",X"44",X"09",
		X"81",X"02",X"00",X"02",X"40",X"C1",X"44",X"09",X"81",X"01",X"02",X"41",X"42",X"C1",X"44",X"09",
		X"81",X"41",X"02",X"02",X"01",X"C1",X"44",X"09",X"81",X"02",X"ED",X"01",X"42",X"C1",X"44",X"09",
		X"81",X"02",X"02",X"02",X"41",X"C1",X"44",X"09",X"81",X"40",X"02",X"02",X"40",X"C1",X"44",X"09",
		X"81",X"02",X"41",X"AD",X"02",X"C1",X"44",X"09",X"81",X"01",X"02",X"02",X"41",X"C1",X"44",X"09",
		X"81",X"02",X"02",X"02",X"42",X"C1",X"44",X"09",X"81",X"ED",X"AD",X"ED",X"AD",X"C1",X"44",X"09",
		X"81",X"02",X"02",X"02",X"42",X"C1",X"44",X"09",X"81",X"02",X"ED",X"01",X"42",X"C1",X"44",X"09",
		X"81",X"02",X"02",X"02",X"02",X"D7",X"44",X"09",X"97",X"02",X"40",X"AD",X"02",X"D9",X"D8",X"44",
		X"07",X"98",X"99",X"41",X"02",X"ED",X"AD",X"DB",X"DA",X"44",X"07",X"9A",X"9B",X"02",X"ED",X"02",
		X"40",X"DE",X"DD",X"44",X"07",X"9D",X"9E",X"ED",X"AD",X"41",X"00",X"E1",X"E0",X"44",X"07",X"A0",
		X"A1",X"42",X"ED",X"01",X"02",X"E4",X"E3",X"44",X"07",X"A3",X"A4",X"02",X"02",X"42",X"ED",X"AD",
		X"E7",X"44",X"07",X"A7",X"41",X"40",X"02",X"AD",X"42",X"42",X"EA",X"44",X"07",X"AA",X"00",X"02",
		X"02",X"02",X"02",X"41",X"D7",X"44",X"07",X"97",X"02",X"02",X"02",X"02",X"02",X"40",X"D9",X"D8",
		X"44",X"05",X"98",X"99",X"ED",X"AD",X"02",X"ED",X"AD",X"02",X"DB",X"DA",X"44",X"05",X"9A",X"9B",
		X"02",X"ED",X"AD",X"AD",X"01",X"02",X"DE",X"DD",X"44",X"05",X"9D",X"9E",X"02",X"02",X"00",X"02",
		X"00",X"01",X"E1",X"E0",X"44",X"05",X"A0",X"A1",X"40",X"01",X"02",X"42",X"ED",X"AD",X"E4",X"E3",
		X"44",X"05",X"A3",X"A4",X"02",X"ED",X"AD",X"AD",X"02",X"ED",X"AD",X"E7",X"44",X"05",X"A7",X"00",
		X"02",X"02",X"ED",X"02",X"02",X"40",X"02",X"EA",X"44",X"05",X"AA",X"02",X"01",X"02",X"02",X"02",
		X"02",X"41",X"42",X"C1",X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",X"02",X"02",X"ED",X"AD",X"C1",
		X"44",X"05",X"81",X"02",X"40",X"42",X"ED",X"ED",X"AD",X"02",X"42",X"C1",X"44",X"05",X"81",X"41",
		X"02",X"ED",X"AD",X"AD",X"42",X"02",X"00",X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"ED",X"ED",
		X"AD",X"42",X"40",X"C1",X"44",X"05",X"81",X"02",X"40",X"42",X"02",X"42",X"ED",X"AD",X"42",X"C1",
		X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",X"AD",X"02",X"02",X"02",X"C1",X"44",X"05",X"81",X"00",
		X"02",X"02",X"ED",X"02",X"02",X"40",X"02",X"C1",X"44",X"05",X"81",X"02",X"01",X"02",X"02",X"02",
		X"02",X"41",X"42",X"C1",X"44",X"05",X"81",X"02",X"42",X"42",X"02",X"01",X"02",X"ED",X"AD",X"C1",
		X"44",X"05",X"81",X"02",X"41",X"42",X"ED",X"02",X"ED",X"AD",X"42",X"C1",X"44",X"05",X"81",X"00",
		X"02",X"ED",X"AD",X"02",X"42",X"02",X"00",X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"42",X"ED",
		X"AD",X"42",X"40",X"C1",X"44",X"05",X"81",X"02",X"40",X"42",X"02",X"AD",X"42",X"42",X"42",X"C1",
		X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",X"41",X"40",X"02",X"02",X"C1",X"44",X"05",X"81",X"ED",
		X"AD",X"02",X"02",X"02",X"02",X"ED",X"AD",X"C1",X"44",X"05",X"81",X"02",X"02",X"ED",X"AD",X"02",
		X"42",X"42",X"02",X"C8",X"C7",X"44",X"04",X"CA",X"77",X"02",X"02",X"02",X"02",X"B4",X"B5",X"02",
		X"6F",X"6E",X"44",X"04",X"7A",X"79",X"F5",X"F4",X"02",X"B5",X"02",X"B4",X"B5",X"71",X"70",X"44",
		X"04",X"7E",X"7F",X"02",X"02",X"02",X"B4",X"B5",X"02",X"02",X"02",X"74",X"73",X"44",X"04",X"C6",
		X"C5",X"B2",X"F2",X"02",X"42",X"42",X"F3",X"F2",X"71",X"70",X"44",X"04",X"C3",X"C2",X"42",X"02",
		X"02",X"B2",X"F2",X"02",X"02",X"02",X"6F",X"6E",X"44",X"04",X"78",X"77",X"B4",X"42",X"42",X"42",
		X"B4",X"B5",X"02",X"71",X"70",X"44",X"04",X"7C",X"79",X"02",X"F5",X"F4",X"02",X"42",X"42",X"02",
		X"02",X"C1",X"44",X"04",X"C3",X"7D",X"02",X"02",X"ED",X"AD",X"42",X"42",X"42",X"42",X"C1",X"44",
		X"05",X"81",X"02",X"02",X"02",X"02",X"ED",X"AD",X"42",X"42",X"C1",X"44",X"05",X"81",X"02",X"AD",
		X"02",X"ED",X"AD",X"02",X"41",X"42",X"C1",X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",X"42",X"42",
		X"42",X"02",X"C1",X"44",X"05",X"81",X"02",X"02",X"ED",X"AD",X"02",X"02",X"40",X"02",X"C1",X"44",
		X"05",X"81",X"02",X"ED",X"AD",X"02",X"ED",X"AD",X"42",X"02",X"C1",X"44",X"05",X"81",X"42",X"AD",
		X"42",X"02",X"02",X"00",X"42",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",X"42",X"ED",X"AD",X"42",
		X"42",X"42",X"C1",X"44",X"05",X"81",X"02",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"C1",X"44",
		X"05",X"81",X"02",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"C1",X"44",X"05",X"81",X"02",X"A8",
		X"E8",X"E8",X"A8",X"E8",X"E8",X"A9",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"42",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"42",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"81",X"02",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"81",X"02",X"9F",X"DF",X"9F",X"DF",X"9F",
		X"9F",X"A2",X"B1",X"44",X"05",X"81",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"C1",X"44",
		X"05",X"81",X"02",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",
		X"02",X"02",X"02",X"B4",X"B5",X"37",X"8A",X"44",X"04",X"96",X"97",X"02",X"F5",X"F4",X"02",X"02",
		X"02",X"02",X"39",X"3A",X"44",X"04",X"2E",X"2F",X"F3",X"02",X"02",X"42",X"F3",X"F2",X"02",X"3F",
		X"3E",X"44",X"04",X"30",X"31",X"42",X"02",X"F3",X"F2",X"02",X"02",X"85",X"86",X"44",X"04",X"33",
		X"34",X"42",X"F5",X"02",X"02",X"F5",X"F4",X"02",X"82",X"83",X"44",X"04",X"30",X"31",X"F5",X"F4",
		X"B4",X"B5",X"42",X"02",X"37",X"38",X"44",X"04",X"2E",X"2F",X"02",X"02",X"42",X"02",X"02",X"02",
		X"02",X"39",X"3C",X"44",X"04",X"30",X"31",X"B2",X"F2",X"42",X"02",X"B4",X"B4",X"B5",X"3D",X"83",
		X"44",X"04",X"81",X"02",X"02",X"42",X"B2",X"02",X"02",X"02",X"37",X"8A",X"44",X"04",X"96",X"97",
		X"42",X"F3",X"F2",X"02",X"F3",X"F2",X"02",X"39",X"3A",X"44",X"04",X"2E",X"2F",X"02",X"02",X"02",
		X"B4",X"02",X"02",X"02",X"3F",X"3E",X"44",X"04",X"30",X"31",X"B4",X"B5",X"02",X"02",X"F5",X"F4",
		X"85",X"86",X"44",X"04",X"33",X"34",X"02",X"42",X"42",X"B2",X"F2",X"B5",X"02",X"82",X"83",X"44",
		X"04",X"30",X"31",X"B4",X"B4",X"B5",X"02",X"02",X"02",X"37",X"38",X"44",X"04",X"2E",X"2F",X"B2",
		X"F2",X"02",X"B4",X"B5",X"02",X"F2",X"39",X"3C",X"44",X"04",X"30",X"31",X"42",X"B4",X"B5",X"02",
		X"B4",X"F4",X"02",X"3D",X"83",X"44",X"04",X"81",X"02",X"B2",X"F2",X"02",X"B2",X"F2",X"02",X"02",
		X"C1",X"44",X"05",X"81",X"02",X"42",X"02",X"02",X"41",X"40",X"02",X"42",X"C1",X"44",X"05",X"81",
		X"02",X"ED",X"AD",X"02",X"42",X"02",X"02",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",X"ED",X"AD",
		X"02",X"02",X"41",X"42",X"C1",X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",X"02",X"02",X"02",X"42",
		X"C1",X"44",X"05",X"81",X"42",X"02",X"42",X"02",X"01",X"02",X"02",X"02",X"C1",X"44",X"05",X"81",
		X"02",X"02",X"02",X"00",X"02",X"ED",X"AD",X"42",X"C1",X"44",X"05",X"81",X"02",X"00",X"42",X"ED",
		X"AD",X"02",X"02",X"02",X"C1",X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",X"02",X"42",X"02",X"02",
		X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"42",X"C1",X"44",X"05",X"81",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"A9",X"B1",X"44",X"05",X"F1",X"E9",X"E8",X"E8",X"E8",
		X"E8",X"E8",X"E8",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",
		X"F0",X"EF",X"06",X"A2",X"B1",X"44",X"05",X"F1",X"E2",X"DF",X"DF",X"DF",X"DF",X"DF",X"DF",X"42",
		X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"C1",X"44",X"05",X"81",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",
		X"BB",X"F8",X"F9",X"F8",X"B9",X"B8",X"FB",X"F0",X"EF",X"06",X"EF",X"0F",X"EF",X"0F",X"EF",X"0F",
		X"EF",X"0F",X"AF",X"FC",X"FE",X"BF",X"BE",X"FF",X"FE",X"BC",X"EF",X"07",X"B0",X"B1",X"44",X"05",
		X"F1",X"F0",X"EF",X"06",X"42",X"C8",X"C7",X"44",X"04",X"CA",X"77",X"42",X"B2",X"F2",X"42",X"02",
		X"02",X"F2",X"6F",X"6E",X"44",X"04",X"7A",X"79",X"42",X"02",X"02",X"B4",X"B4",X"F4",X"42",X"71",
		X"70",X"44",X"04",X"7E",X"7F",X"42",X"B4",X"B5",X"42",X"42",X"B4",X"B5",X"42",X"74",X"73",X"44",
		X"04",X"C6",X"C5",X"42",X"42",X"B2",X"F2",X"02",X"F5",X"F4",X"71",X"70",X"44",X"04",X"C3",X"C2",
		X"42",X"F3",X"F2",X"42",X"42",X"F4",X"42",X"42",X"6F",X"6E",X"44",X"04",X"78",X"77",X"42",X"42",
		X"B2",X"F2",X"42",X"B2",X"F2",X"71",X"70",X"44",X"04",X"7C",X"79",X"F5",X"B4",X"B5",X"42",X"B2",
		X"F2",X"42",X"42",X"C1",X"44",X"04",X"C3",X"7D",X"B2",X"F2",X"42",X"42",X"02",X"02",X"02",X"02",
		X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"C1",X"44",X"05",X"81",
		X"42",X"42",X"42",X"42",X"E8",X"E8",X"E8",X"A9",X"B1",X"44",X"05",X"F1",X"E9",X"E8",X"E8",X"E8",
		X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",
		X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",
		X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",
		X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",
		X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",
		X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",
		X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",
		X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",
		X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",
		X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",
		X"EF",X"03",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"03",X"EF",X"03",X"B0",X"B1",X"44",X"05",
		X"F1",X"F0",X"EF",X"03",X"9F",X"9F",X"9F",X"A2",X"B1",X"44",X"05",X"F1",X"E2",X"9F",X"9F",X"9F",
		X"42",X"42",X"42",X"42",X"C1",X"44",X"05",X"81",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"42",
		X"C1",X"44",X"05",X"81",X"42",X"42",X"42",X"42",X"02",X"41",X"42",X"42",X"66",X"44",X"05",X"26",
		X"02",X"02",X"02",X"02",X"02",X"02",X"40",X"48",X"47",X"44",X"05",X"07",X"08",X"ED",X"AD",X"02",
		X"02",X"ED",X"AD",X"4E",X"4D",X"44",X"05",X"0D",X"0E",X"02",X"ED",X"AD",X"02",X"00",X"42",X"53",
		X"52",X"44",X"05",X"12",X"13",X"02",X"02",X"ED",X"AD",X"02",X"42",X"66",X"44",X"07",X"26",X"01",
		X"02",X"02",X"ED",X"AD",X"48",X"47",X"44",X"07",X"07",X"08",X"ED",X"AD",X"AD",X"02",X"4E",X"4D",
		X"44",X"07",X"0D",X"0E",X"00",X"02",X"02",X"42",X"53",X"52",X"44",X"07",X"12",X"13",X"02",X"02",
		X"02",X"02",X"66",X"44",X"09",X"26",X"02",X"02",X"01",X"48",X"47",X"44",X"09",X"07",X"08",X"02",
		X"02",X"4E",X"4D",X"44",X"09",X"0D",X"0E",X"ED",X"AD",X"53",X"52",X"44",X"09",X"12",X"13",X"00",
		X"02",X"66",X"44",X"04",X"96",X"A6",X"D6",X"44",X"04",X"26",X"02",X"48",X"47",X"44",X"04",X"2E",
		X"8B",X"6E",X"44",X"04",X"07",X"08",X"4E",X"4D",X"44",X"04",X"A0",X"8B",X"E0",X"44",X"04",X"0D",
		X"0E",X"53",X"52",X"44",X"04",X"A3",X"8B",X"E3",X"44",X"04",X"12",X"13",X"C1",X"44",X"05",X"81",
		X"00",X"C1",X"44",X"05",X"81",X"C1",X"44",X"05",X"81",X"41",X"C1",X"44",X"05",X"81",X"C1",X"44",
		X"05",X"81",X"40",X"C1",X"44",X"05",X"81",X"C1",X"44",X"05",X"81",X"01",X"C1",X"44",X"05",X"81",
		X"C1",X"44",X"05",X"81",X"00",X"C1",X"44",X"05",X"81",X"C1",X"44",X"05",X"81",X"41",X"C1",X"44",
		X"05",X"81",X"C1",X"44",X"05",X"81",X"40",X"C1",X"44",X"05",X"81",X"C1",X"44",X"05",X"81",X"01",
		X"C1",X"44",X"05",X"81",X"C1",X"44",X"05",X"97",X"00",X"D7",X"44",X"05",X"81",X"C1",X"44",X"04",
		X"98",X"99",X"41",X"D9",X"D8",X"44",X"04",X"81",X"C1",X"44",X"04",X"9A",X"9B",X"40",X"DB",X"DA",
		X"44",X"04",X"81",X"C1",X"44",X"04",X"9D",X"9E",X"41",X"DE",X"DD",X"44",X"04",X"81",X"C1",X"44",
		X"04",X"A0",X"A1",X"00",X"E1",X"E0",X"44",X"04",X"81",X"C1",X"44",X"04",X"A3",X"A4",X"01",X"E4",
		X"E3",X"44",X"04",X"81",X"C1",X"44",X"04",X"A7",X"02",X"40",X"42",X"E7",X"44",X"04",X"81",X"C1",
		X"44",X"04",X"AA",X"01",X"02",X"41",X"EA",X"44",X"04",X"81",X"C1",X"44",X"04",X"81",X"02",X"02",
		X"02",X"EA",X"44",X"04",X"81",X"B1",X"44",X"04",X"F1",X"E9",X"A8",X"A9",X"B1",X"44",X"04",X"F1",
		X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",
		X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",
		X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",
		X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",
		X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",
		X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",
		X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",
		X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",
		X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",
		X"44",X"04",X"F1",X"F0",X"AF",X"B0",X"B1",X"44",X"04",X"F1",X"B1",X"44",X"04",X"F1",X"E2",X"DF",
		X"A2",X"B1",X"44",X"04",X"F1",X"C1",X"44",X"04",X"81",X"02",X"02",X"02",X"C1",X"44",X"04",X"81",
		X"C1",X"44",X"04",X"26",X"02",X"40",X"42",X"66",X"44",X"04",X"81",X"C1",X"44",X"04",X"07",X"08",
		X"01",X"48",X"47",X"44",X"04",X"81",X"C1",X"44",X"04",X"0D",X"0E",X"00",X"4E",X"4D",X"44",X"04",
		X"81",X"C1",X"44",X"04",X"12",X"13",X"41",X"53",X"52",X"44",X"04",X"81",X"C1",X"44",X"05",X"81",
		X"40",X"C1",X"44",X"05",X"81",X"C1",X"44",X"05",X"81",X"01",X"C1",X"44",X"05",X"81",X"C1",X"44",
		X"05",X"81",X"00",X"C1",X"44",X"05",X"81",X"C1",X"44",X"05",X"81",X"41",X"C1",X"44",X"05",X"81",
		X"D7",X"44",X"05",X"81",X"40",X"C1",X"44",X"05",X"97",X"D9",X"D8",X"44",X"04",X"81",X"01",X"C1",
		X"44",X"04",X"98",X"99",X"DB",X"DA",X"44",X"04",X"81",X"00",X"C1",X"44",X"04",X"9A",X"9B",X"DE",
		X"DD",X"44",X"04",X"78",X"5C",X"38",X"44",X"04",X"9D",X"9E",X"E1",X"E0",X"44",X"04",X"1A",X"1C",
		X"5A",X"44",X"04",X"A0",X"A1",X"E4",X"E3",X"44",X"04",X"1A",X"1C",X"5A",X"44",X"04",X"A3",X"A4",
		X"02",X"66",X"44",X"04",X"05",X"1C",X"5A",X"44",X"04",X"81",X"02",X"39",X"3A",X"44",X"03",X"24",
		X"25",X"22",X"23",X"44",X"03",X"33",X"34",X"01",X"3F",X"3E",X"44",X"03",X"2A",X"2B",X"28",X"44",
		X"04",X"30",X"31",X"ED",X"86",X"44",X"04",X"05",X"06",X"03",X"44",X"04",X"81",X"ED",X"AD",X"83",
		X"44",X"03",X"0B",X"0C",X"09",X"0A",X"44",X"04",X"81",X"02",X"02",X"44",X"04",X"10",X"11",X"0F",
		X"44",X"05",X"81",X"02",X"ED",X"44",X"03",X"0B",X"0C",X"09",X"0A",X"44",X"05",X"81",X"ED",X"AD",
		X"44",X"03",X"10",X"11",X"0F",X"44",X"06",X"81",X"02",X"02",X"04",X"04",X"0B",X"0C",X"09",X"0A",
		X"44",X"06",X"81",X"02",X"02",X"04",X"04",X"10",X"11",X"0F",X"44",X"07",X"81",X"41",X"00",X"04",
		X"0B",X"0C",X"09",X"0A",X"44",X"07",X"81",X"02",X"ED",X"04",X"10",X"11",X"0F",X"44",X"08",X"81",
		X"02",X"ED",X"0B",X"0C",X"09",X"0A",X"44",X"08",X"81",X"40",X"02",X"10",X"8D",X"28",X"44",X"09",
		X"81",X"02",X"02",X"0C",X"92",X"70",X"44",X"09",X"81",X"ED",X"AD",X"94",X"42",X"C1",X"44",X"09",
		X"81",X"42",X"42",X"42",X"C1",X"44",X"04",X"1A",X"1C",X"45",X"44",X"04",X"26",X"02",X"AD",X"74",
		X"73",X"44",X"03",X"63",X"62",X"65",X"64",X"44",X"03",X"7A",X"79",X"02",X"71",X"70",X"44",X"04",
		X"68",X"6B",X"6A",X"44",X"03",X"7E",X"7F",X"41",X"42",X"C1",X"44",X"04",X"43",X"46",X"45",X"44",
		X"04",X"C6",X"42",X"40",X"C1",X"44",X"04",X"4A",X"49",X"4C",X"4B",X"44",X"03",X"C3",X"ED",X"AD",
		X"C1",X"44",X"05",X"4F",X"51",X"50",X"44",X"04",X"AD",X"42",X"C1",X"44",X"05",X"4A",X"49",X"4C",
		X"4B",X"44",X"03",X"02",X"02",X"C1",X"44",X"06",X"4F",X"51",X"50",X"44",X"03",X"42",X"42",X"C1",
		X"44",X"06",X"4A",X"49",X"4C",X"4B",X"04",X"04",X"ED",X"AD",X"C1",X"44",X"07",X"4F",X"51",X"50",
		X"04",X"04",X"40",X"42",X"C1",X"44",X"07",X"4A",X"49",X"4C",X"4B",X"04",X"AD",X"42",X"C1",X"44",
		X"08",X"4F",X"51",X"50",X"04",X"02",X"02",X"C1",X"44",X"08",X"4A",X"49",X"4C",X"4B",X"01",X"00",
		X"C1",X"44",X"09",X"68",X"CD",X"50",X"AD",X"42",X"C1",X"44",X"09",X"30",X"D2",X"4C",X"02",X"02",
		X"C1",X"44",X"09",X"81",X"01",X"D4",X"42",X"C1",X"44",X"05",X"CA",X"77",X"42",X"02",X"42",X"42",
		X"42",X"02",X"42",X"C1",X"44",X"05",X"7A",X"79",X"00",X"02",X"ED",X"AD",X"42",X"02",X"02",X"C1",
		X"44",X"05",X"7E",X"7F",X"42",X"42",X"02",X"02",X"ED",X"AD",X"02",X"C1",X"44",X"06",X"C6",X"C5",
		X"41",X"42",X"42",X"42",X"02",X"42",X"C1",X"44",X"06",X"C3",X"C2",X"42",X"42",X"ED",X"AD",X"02",
		X"42",X"C1",X"44",X"07",X"78",X"77",X"00",X"42",X"42",X"ED",X"02",X"C1",X"44",X"07",X"7C",X"79",
		X"42",X"41",X"42",X"02",X"02",X"C1",X"44",X"07",X"C3",X"7D",X"42",X"42",X"ED",X"AD",X"42",X"C1",
		X"44",X"08",X"CA",X"77",X"42",X"42",X"02",X"42",X"C1",X"44",X"08",X"7A",X"79",X"ED",X"AD",X"02",
		X"02",X"C1",X"44",X"08",X"7E",X"7F",X"42",X"42",X"40",X"02",X"C1",X"44",X"05",X"96",X"E6",X"D6",
		X"04",X"C6",X"C5",X"41",X"02",X"42",X"C1",X"44",X"05",X"2E",X"CB",X"6E",X"04",X"C3",X"C2",X"42",
		X"ED",X"42",X"C1",X"44",X"05",X"A3",X"CD",X"E3",X"04",X"04",X"78",X"77",X"02",X"02",X"C1",X"44",
		X"05",X"81",X"D2",X"70",X"04",X"04",X"7C",X"79",X"41",X"02",X"C1",X"44",X"05",X"81",X"42",X"74",
		X"73",X"04",X"C3",X"7D",X"02",X"02",X"C1",X"44",X"05",X"81",X"41",X"E4",X"E3",X"04",X"04",X"81",
		X"02",X"42",X"C1",X"44",X"05",X"81",X"42",X"40",X"E7",X"04",X"04",X"81",X"02",X"02",X"C1",X"44",
		X"05",X"81",X"01",X"42",X"EA",X"04",X"04",X"81",X"02",X"02",X"C1",X"44",X"05",X"81",X"02",X"00",
		X"D7",X"04",X"04",X"81",X"02",X"42",X"C1",X"44",X"05",X"81",X"41",X"02",X"D9",X"D8",X"04",X"81",
		X"02",X"42",X"C1",X"44",X"05",X"81",X"42",X"01",X"DB",X"DA",X"04",X"81",X"02",X"42",X"C1",X"44",
		X"05",X"81",X"40",X"02",X"DE",X"DD",X"04",X"81",X"02",X"42",X"C1",X"44",X"05",X"81",X"02",X"00",
		X"E1",X"E0",X"04",X"81",X"42",X"02",X"C1",X"44",X"05",X"81",X"02",X"01",X"E4",X"E3",X"04",X"81",
		X"02",X"42",X"C1",X"44",X"05",X"81",X"42",X"00",X"42",X"66",X"04",X"26",X"02",X"02",X"C1",X"44",
		X"05",X"81",X"42",X"41",X"48",X"47",X"04",X"07",X"08",X"A9",X"B1",X"44",X"05",X"F1",X"E9",X"E8",
		X"E5",X"67",X"AF",X"27",X"A5",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",X"05",X"F1",X"F0",X"EF",X"06",X"B0",X"B1",X"44",
		X"05",X"F1",X"F0",X"EF",X"06",X"A2",X"B1",X"44",X"05",X"F1",X"E2",X"EE",X"72",X"EF",X"04",X"42",
		X"C1",X"44",X"05",X"81",X"02",X"02",X"D3",X"D0",X"EF",X"03",X"02",X"C1",X"44",X"05",X"81",X"02",
		X"02",X"C0",X"7B",X"EF",X"03",X"02",X"C1",X"44",X"05",X"81",X"02",X"41",X"69",X"5B",X"EF",X"03",
		X"42",X"C1",X"44",X"05",X"81",X"02",X"42",X"6F",X"5B",X"EF",X"03",X"42",X"C1",X"44",X"05",X"81",
		X"02",X"40",X"42",X"D3",X"D0",X"AF",X"AF",X"42",X"C1",X"44",X"05",X"81",X"41",X"42",X"42",X"69",
		X"5B",X"AF",X"AF",X"42",X"C1",X"44",X"05",X"81",X"42",X"02",X"42",X"6F",X"7B",X"AF",X"AF",X"02",
		X"C1",X"44",X"05",X"81",X"42",X"ED",X"AD",X"02",X"D3",X"72",X"AF",X"42",X"C1",X"44",X"05",X"81",
		X"02",X"02",X"42",X"01",X"69",X"5B",X"AF",X"02",X"C1",X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",
		X"C0",X"5B",X"AF",X"02",X"C1",X"44",X"05",X"81",X"02",X"02",X"42",X"42",X"69",X"7B",X"AF",X"42",
		X"C1",X"44",X"05",X"81",X"02",X"42",X"42",X"01",X"6F",X"5B",X"AF",X"42",X"C1",X"44",X"05",X"81",
		X"02",X"40",X"42",X"42",X"42",X"D3",X"D0",X"42",X"C1",X"44",X"05",X"81",X"41",X"42",X"42",X"ED",
		X"AD",X"39",X"5B",X"42",X"C1",X"44",X"05",X"81",X"42",X"02",X"42",X"42",X"42",X"6F",X"7B",X"02",
		X"C1",X"44",X"05",X"81",X"42",X"ED",X"AD",X"02",X"42",X"42",X"D3",X"42",X"C1",X"44",X"05",X"81",
		X"02",X"02",X"42",X"02",X"01",X"42",X"6F",X"02",X"C1",X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",
		X"42",X"42",X"02",X"02",X"42",X"C0",X"7B",X"EF",X"07",X"1B",X"29",X"59",X"58",X"02",X"42",X"C0",
		X"7B",X"EF",X"07",X"1B",X"29",X"59",X"58",X"02",X"42",X"69",X"5B",X"EF",X"07",X"3B",X"29",X"59",
		X"1F",X"02",X"42",X"C9",X"C4",X"EF",X"07",X"1B",X"29",X"6C",X"5F",X"A8",X"E5",X"67",X"EF",X"08",
		X"84",X"29",X"59",X"58",X"EF",X"0B",X"90",X"29",X"5E",X"5D",X"EF",X"0B",X"3B",X"80",X"59",X"58",
		X"EF",X"0B",X"1B",X"29",X"6C",X"1F",X"EF",X"0B",X"1B",X"29",X"59",X"58",X"EF",X"0B",X"3B",X"80",
		X"59",X"1F",X"EF",X"0B",X"1B",X"29",X"6C",X"5F",X"EF",X"0B",X"84",X"29",X"59",X"58",X"EF",X"0B",
		X"90",X"29",X"5E",X"5D",X"EF",X"0B",X"3B",X"80",X"59",X"58",X"EF",X"0B",X"1B",X"29",X"6C",X"1F",
		X"EF",X"0B",X"1B",X"29",X"59",X"58",X"72",X"EF",X"0A",X"3B",X"80",X"5E",X"5F",X"5B",X"EF",X"0A",
		X"1B",X"29",X"5F",X"58",X"D3",X"D0",X"EF",X"09",X"84",X"29",X"1F",X"5F",X"C0",X"5B",X"EF",X"09",
		X"90",X"80",X"6C",X"58",X"5F",X"D3",X"72",X"EF",X"08",X"1B",X"29",X"76",X"5F",X"18",X"5F",X"D3",
		X"D0",X"EF",X"07",X"1B",X"29",X"5F",X"5D",X"8E",X"2C",X"39",X"7B",X"EF",X"07",X"3B",X"80",X"59",
		X"5D",X"42",X"42",X"69",X"5B",X"EF",X"07",X"1B",X"29",X"5E",X"5D",X"35",X"36",X"C0",X"7B",X"EF",
		X"07",X"3B",X"80",X"5E",X"5F",X"1D",X"19",X"69",X"5B",X"EF",X"07",X"1B",X"29",X"59",X"58",X"18",
		X"35",X"36",X"D3",X"D0",X"EF",X"06",X"84",X"29",X"5E",X"5F",X"42",X"18",X"19",X"C0",X"7B",X"EF",
		X"06",X"90",X"80",X"6C",X"58",X"42",X"1D",X"1E",X"69",X"C4",X"EF",X"06",X"1B",X"29",X"76",X"75",
		X"18",X"18",X"19",X"C0",X"7B",X"EF",X"06",X"1B",X"29",X"59",X"5D",X"8E",X"2C",X"2D",X"69",X"5B",
		X"EF",X"06",X"3B",X"80",X"59",X"5D",X"AB",X"35",X"36",X"69",X"5B",X"EF",X"06",X"1B",X"29",X"5E",
		X"5D",X"1F",X"1D",X"1E",X"69",X"5B",X"EF",X"06",X"3B",X"80",X"6D",X"6C",X"1D",X"2C",X"2D",X"69",
		X"C4",X"EF",X"06",X"1B",X"29",X"76",X"75",X"5F",X"35",X"42",X"6F",X"D0",X"EF",X"06",X"84",X"29",
		X"59",X"6C",X"1F",X"2D",X"02",X"85",X"7B",X"EF",X"06",X"90",X"80",X"59",X"1F",X"1F",X"AB",X"35",
		X"69",X"C4",X"EF",X"06",X"3B",X"29",X"5E",X"5D",X"18",X"18",X"19",X"C0",X"D0",X"EF",X"06",X"1B",
		X"29",X"59",X"5D",X"18",X"18",X"19",X"69",X"5B",X"EF",X"06",X"3B",X"80",X"6D",X"6C",X"1F",X"18",
		X"1E",X"69",X"5B",X"EF",X"06",X"1B",X"29",X"76",X"75",X"1F",X"1D",X"1E",X"69",X"5B",X"EF",X"06",
		X"3B",X"80",X"5E",X"5D",X"1D",X"1D",X"1E",X"C0",X"7B",X"EF",X"06",X"1B",X"29",X"59",X"58",X"18",
		X"6C",X"19",X"69",X"5B",X"EF",X"06",X"84",X"29",X"6D",X"6C",X"1F",X"1F",X"19",X"C0",X"7B",X"AF",
		X"AF",X"3B",X"D0",X"AF",X"AF",X"90",X"80",X"42",X"42",X"42",X"75",X"1E",X"69",X"5B",X"AF",X"AF",
		X"1B",X"7B",X"AF",X"AF",X"1B",X"29",X"76",X"75",X"18",X"19",X"2D",X"C9",X"C4",X"AF",X"AF",X"84",
		X"5B",X"AF",X"AF",X"1B",X"29",X"59",X"5D",X"18",X"1E",X"39",X"7B",X"EF",X"07",X"3B",X"80",X"5E",
		X"5F",X"18",X"19",X"69",X"5B",X"EF",X"07",X"1B",X"29",X"59",X"58",X"02",X"1E",X"C0",X"7B",X"EF",
		X"07",X"3B",X"80",X"5E",X"5F",X"1D",X"19",X"69",X"5B",X"EF",X"07",X"1B",X"29",X"59",X"58",X"18",
		X"35",X"36",X"D3",X"D0",X"EF",X"06",X"84",X"29",X"5E",X"5F",X"42",X"18",X"19",X"C0",X"7B",X"EF",
		X"06",X"90",X"80",X"6C",X"58",X"42",X"1D",X"1E",X"69",X"5B",X"EF",X"06",X"1B",X"29",X"76",X"75",
		X"18",X"18",X"2D",X"C9",X"C4",X"EF",X"06",X"1B",X"29",X"59",X"5D",X"8E",X"2C",X"39",X"7B",X"EF",
		X"07",X"3B",X"80",X"59",X"5D",X"AB",X"35",X"69",X"5B",X"EF",X"07",X"1B",X"29",X"5E",X"5D",X"02",
		X"1E",X"C0",X"7B",X"EF",X"07",X"84",X"89",X"6D",X"18",X"1D",X"19",X"69",X"5B",X"EF",X"03",X"32",
		X"AE",X"72",X"AF",X"AF",X"27",X"A5",X"A8",X"18",X"35",X"36",X"D3",X"D0",X"AF",X"AF",X"3B",X"93",
		X"D3",X"D0",X"AF",X"AF",X"AF",X"32",X"42",X"18",X"19",X"C0",X"7B",X"AF",X"AF",X"1B",X"79",X"C9",
		X"C4",X"AF",X"AF",X"90",X"93",X"42",X"1D",X"1E",X"69",X"C4",X"AF",X"AF",X"27",X"E5",X"67",X"AF",
		X"AF",X"AF",X"1B",X"9B",X"18",X"18",X"19",X"C0",X"7B",X"EF",X"06",X"32",X"AE",X"93",X"02",X"8E",
		X"2C",X"2D",X"69",X"5B",X"EF",X"06",X"1B",X"34",X"76",X"75",X"AB",X"35",X"36",X"69",X"5B",X"EF",
		X"06",X"1B",X"29",X"5E",X"5D",X"8E",X"2C",X"2D",X"6F",X"5B",X"EF",X"06",X"3B",X"80",X"5E",X"5D",
		X"A5",X"89",X"02",X"42",X"D3",X"EE",X"72",X"EF",X"04",X"1B",X"29",X"59",X"58",X"AF",X"84",X"E5",
		X"A5",X"89",X"D3",X"D0",X"EF",X"04",X"84",X"29",X"6D",X"6C",X"EF",X"04",X"84",X"E5",X"67",X"EF",
		X"04",X"90",X"80",X"76",X"75",X"EF",X"0B",X"1B",X"29",X"6D",X"6C",X"DF",X"EE",X"72",X"EF",X"08",
		X"1B",X"29",X"76",X"75",X"AB",X"35",X"D3",X"D0",X"EF",X"07",X"3B",X"80",X"5E",X"5F",X"42",X"18",
		X"69",X"5B",X"EF",X"07",X"1B",X"29",X"59",X"58",X"5F",X"C0",X"7B",X"EF",X"0A",X"3B",X"A4",X"1D",
		X"4E",X"5B",X"EF",X"04",X"3B",X"D0",X"EF",X"04",X"1B",X"A4",X"18",X"C0",X"7B",X"EF",X"03",X"90",
		X"93",X"D3",X"72",X"EF",X"03",X"1B",X"A4",X"1D",X"69",X"C4",X"EF",X"03",X"1B",X"A4",X"6F",X"7B",
		X"EF",X"03",X"3B",X"A4",X"5F",X"69",X"D0",X"EF",X"03",X"3B",X"A4",X"48",X"5B",X"EF",X"03",X"1B",
		X"A4",X"18",X"C0",X"7B",X"AF",X"AF",X"32",X"93",X"02",X"C9",X"C4",X"EF",X"03",X"3B",X"A4",X"1D",
		X"69",X"5B",X"AF",X"AF",X"1B",X"2F",X"85",X"C4",X"EF",X"03",X"32",X"93",X"02",X"1F",X"69",X"5B",
		X"AF",X"AF",X"3B",X"A4",X"69",X"D0",X"EF",X"03",X"1B",X"2F",X"02",X"5F",X"C0",X"5B",X"AF",X"AF",
		X"1B",X"A4",X"C9",X"C4",X"EF",X"03",X"1B",X"29",X"02",X"58",X"39",X"5B",X"AF",X"32",X"93",X"39",
		X"C4",X"EF",X"04",X"3B",X"2F",X"5F",X"42",X"C0",X"7B",X"AF",X"3B",X"2F",X"6F",X"D0",X"EF",X"04",
		X"1B",X"79",X"6C",X"42",X"71",X"70",X"04",X"30",X"31",X"39",X"7B",X"EF",X"04",X"84",X"0E",X"42",
		X"01",X"42",X"C1",X"04",X"81",X"02",X"69",X"5B",X"EF",X"04",X"90",X"2F",X"75",X"42",X"42",X"66",
		X"04",X"97",X"42",X"C0",X"C4",X"EF",X"04",X"1B",X"A4",X"5F",X"00",X"48",X"47",X"98",X"99",X"42",
		X"69",X"D0",X"EF",X"04",X"3B",X"79",X"1F",X"42",X"4E",X"4D",X"9A",X"9B",X"42",X"C0",X"5B",X"EF",
		X"04",X"1B",X"29",X"58",X"42",X"53",X"52",X"9D",X"9E",X"02",X"69",X"7B",X"EF",X"04",X"1B",X"29",
		X"02",X"42",X"66",X"04",X"A0",X"A1",X"02",X"69",X"5B",X"EF",X"04",X"3B",X"2F",X"5F",X"48",X"47",
		X"04",X"30",X"31",X"42",X"C0",X"5B",X"EF",X"04",X"1B",X"79",X"6C",X"3F",X"3E",X"33",X"34",X"42",
		X"42",X"69",X"7B",X"EF",X"04",X"84",X"0E",X"42",X"86",X"04",X"30",X"31",X"42",X"42",X"69",X"5B",
		X"EF",X"04",X"90",X"2F",X"75",X"83",X"33",X"34",X"42",X"42",X"42",X"C0",X"C4",X"EF",X"04",X"1B",
		X"A4",X"5F",X"04",X"30",X"31",X"75",X"35",X"36",X"69",X"D0",X"EF",X"04",X"3B",X"79",X"1F",X"33",
		X"34",X"02",X"59",X"5F",X"1E",X"C0",X"5B",X"EF",X"04",X"1B",X"29",X"58",X"30",X"31",X"75",X"1F",
		X"5F",X"2D",X"C9",X"C4",X"EF",X"04",X"1B",X"29",X"58",X"34",X"76",X"5F",X"1D",X"2D",X"39",X"5B",
		X"EF",X"05",X"3B",X"2F",X"6C",X"31",X"59",X"1F",X"19",X"02",X"C9",X"C4",X"EF",X"05",X"84",X"79",
		X"02",X"02",X"1F",X"1F",X"19",X"85",X"C4",X"EF",X"06",X"90",X"2F",X"75",X"02",X"1F",X"1F",X"2D",
		X"69",X"D0",X"EF",X"06",X"1B",X"A1",X"18",X"02",X"1D",X"19",X"02",X"C0",X"7B",X"EF",X"06",X"3B",
		X"A1",X"59",X"02",X"1D",X"18",X"35",X"69",X"5B",X"EF",X"06",X"1B",X"79",X"02",X"5F",X"5F",X"1D",
		X"2C",X"C9",X"C4",X"EF",X"06",X"3B",X"2F",X"1F",X"18",X"1F",X"58",X"39",X"5B",X"EF",X"07",X"1B",
		X"29",X"58",X"02",X"5F",X"58",X"6F",X"D0",X"EF",X"07",X"1B",X"2F",X"6C",X"1D",X"18",X"19",X"85",
		X"5B",X"EF",X"07",X"84",X"79",X"18",X"5F",X"1F",X"1F",X"C0",X"7B",X"EF",X"07",X"90",X"2F",X"75",
		X"02",X"1F",X"19",X"39",X"C4",X"EF",X"07",X"1B",X"A1",X"18",X"5F",X"1D",X"5F",X"69",X"5B",X"EF",
		X"07",X"3B",X"A1",X"59",X"02",X"1D",X"1E",X"39",X"7B",X"EF",X"07",X"1B",X"79",X"18",X"5F",X"5F",
		X"5D",X"6F",X"5B",X"EF",X"07",X"3B",X"2F",X"58",X"18",X"1F",X"58",X"39",X"5B",X"EF",X"07",X"84",
		X"29",X"58",X"02",X"18",X"5F",X"6F",X"D0",X"EF",X"07",X"90",X"2F",X"6C",X"1D",X"18",X"2C",X"85",
		X"5B",X"EF",X"03",X"32",X"D0",X"AF",X"AF",X"1B",X"79",X"18",X"5F",X"1F",X"42",X"C9",X"C4",X"EF",
		X"03",X"84",X"67",X"AF",X"AF",X"1B",X"2F",X"75",X"02",X"19",X"E4",X"7B",X"EF",X"08",X"84",X"A1",
		X"18",X"5F",X"58",X"85",X"5B",X"AF",X"AF",X"90",X"7B",X"EF",X"04",X"90",X"A1",X"59",X"02",X"5F",
		X"69",X"C4",X"AF",X"AF",X"27",X"67",X"EF",X"04",X"1B",X"79",X"18",X"5F",X"5F",X"69",X"5B",X"EF",
		X"08",X"1B",X"2F",X"58",X"18",X"5F",X"C0",X"7B",X"EF",X"08",X"84",X"29",X"58",X"02",X"18",X"6F",
		X"5B",X"EF",X"08",X"90",X"2F",X"6C",X"1D",X"18",X"39",X"5B",X"EF",X"08",X"1B",X"79",X"18",X"5F",
		X"1F",X"69",X"D0",X"EF",X"08",X"1B",X"2F",X"75",X"02",X"19",X"E4",X"7B",X"EF",X"08",X"84",X"A1",
		X"18",X"5F",X"58",X"85",X"5B",X"EF",X"08",X"90",X"A1",X"59",X"02",X"5F",X"69",X"C4",X"EF",X"08",
		X"1B",X"79",X"18",X"5F",X"5F",X"69",X"5B",X"EF",X"08",X"1B",X"2F",X"58",X"18",X"5F",X"C0",X"7B",
		X"EF",X"08",X"84",X"29",X"58",X"1F",X"58",X"6F",X"5B",X"EF",X"08",X"90",X"2F",X"6C",X"1D",X"02",
		X"C9",X"67",X"EF",X"08",X"1B",X"79",X"18",X"5F",X"E4",X"7B",X"EF",X"09",X"1B",X"2F",X"75",X"19",
		X"85",X"5B",X"EF",X"09",X"84",X"A1",X"18",X"5F",X"DB",X"C4",X"EF",X"09",X"90",X"A1",X"59",X"5F",
		X"E1",X"5B",X"EF",X"09",X"1B",X"79",X"18",X"5F",X"39",X"7B",X"EF",X"09",X"1B",X"2F",X"58",X"18",
		X"69",X"5B",X"EF",X"09",X"1B",X"29",X"58",X"1F",X"6F",X"D0",X"EF",X"09",X"3B",X"2F",X"6C",X"1D",
		X"E4",X"5B",X"EF",X"09",X"1B",X"79",X"18",X"5F",X"E4",X"7B",X"EF",X"09",X"1B",X"2F",X"75",X"19",
		X"85",X"5B",X"EF",X"09",X"84",X"A1",X"18",X"5F",X"DB",X"C4",X"EF",X"09",X"90",X"A1",X"59",X"5F",
		X"E1",X"5B",X"EF",X"09",X"1B",X"79",X"18",X"5F",X"39",X"7B",X"EF",X"09",X"1B",X"2F",X"58",X"18",
		X"5F",X"C0",X"7B",X"EF",X"07",X"1B",X"80",X"5F",X"1F",X"02",X"18",X"6F",X"5B",X"EF",X"07",X"3B",
		X"2F",X"59",X"5F",X"1D",X"18",X"39",X"C4",X"EF",X"07",X"84",X"89",X"6C",X"5F",X"5F",X"1F",X"69",
		X"D0",X"EF",X"08",X"1B",X"A4",X"18",X"02",X"19",X"E4",X"7B",X"EF",X"08",X"84",X"A1",X"18",X"5F",
		X"58",X"85",X"5B",X"EF",X"08",X"90",X"A1",X"59",X"02",X"5F",X"69",X"5B",X"EF",X"08",X"1B",X"79",
		X"18",X"5F",X"5F",X"69",X"5B",X"EF",X"08",X"1B",X"2F",X"58",X"18",X"69",X"5B",X"EF",X"09",X"1B",
		X"29",X"58",X"1F",X"6F",X"D0",X"EF",X"04",X"3B",X"D0",X"AF",X"AF",X"AF",X"3B",X"2F",X"6C",X"58",
		X"E4",X"5B",X"EF",X"04",X"1B",X"C4",X"AF",X"AF",X"90",X"93",X"75",X"18",X"19",X"E4",X"7B",X"EF",
		X"04",X"84",X"D0",X"AF",X"AF",X"1B",X"2F",X"1F",X"18",X"58",X"35",X"D3",X"D0",X"EF",X"07",X"3B",
		X"79",X"1F",X"18",X"5F",X"58",X"DB",X"C4",X"EF",X"07",X"1B",X"80",X"59",X"1F",X"5F",X"5F",X"E1",
		X"5B",X"AF",X"AF",X"90",X"72",X"EF",X"03",X"84",X"29",X"18",X"18",X"5F",X"1E",X"39",X"7B",X"AF",
		X"AF",X"1B",X"D0",X"EF",X"03",X"90",X"80",X"5F",X"58",X"18",X"5F",X"C0",X"7B",X"EF",X"08",X"84",
		X"89",X"58",X"1F",X"58",X"6F",X"5B",X"EF",X"09",X"1B",X"79",X"1D",X"02",X"C9",X"67",X"EF",X"09",
		X"1B",X"2F",X"5F",X"E4",X"7B",X"EF",X"0A",X"84",X"29",X"19",X"85",X"5B",X"EF",X"0A",X"90",X"2F",
		X"5F",X"DB",X"C4",X"EF",X"0A",X"3B",X"79",X"5F",X"E1",X"5B",X"EF",X"0A",X"1B",X"2F",X"5F",X"39",
		X"7B",X"EF",X"0A",X"3B",X"A4",X"18",X"69",X"5B",X"EF",X"0A",X"1B",X"29",X"1F",X"6F",X"D0",X"EF",
		X"0A",X"3B",X"2F",X"1D",X"E4",X"5B",X"EF",X"0A",X"1B",X"79",X"5F",X"E4",X"7B",X"EF",X"0A",X"1B",
		X"2F",X"19",X"85",X"5B",X"EF",X"0A",X"84",X"A1",X"5F",X"DB",X"C4",X"EF",X"0A",X"90",X"A1",X"5F",
		X"E1",X"5B",X"EF",X"0A",X"1B",X"79",X"5F",X"39",X"7B",X"EF",X"0A",X"1B",X"2F",X"02",X"C1",X"44",
		X"05",X"81",X"02",X"40",X"02",X"02",X"02",X"02",X"02",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",
		X"42",X"ED",X"AD",X"02",X"02",X"42",X"C1",X"44",X"05",X"81",X"02",X"41",X"02",X"02",X"02",X"02",
		X"02",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"40",X"02",X"02",X"02",X"42",X"C1",X"44",
		X"05",X"81",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"C1",X"44",X"05",X"81",X"02",X"00",
		X"02",X"02",X"02",X"ED",X"AD",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"02",X"02",X"02",
		X"37",X"02",X"C1",X"44",X"05",X"81",X"02",X"ED",X"AD",X"02",X"02",X"02",X"3F",X"02",X"C1",X"44",
		X"05",X"81",X"02",X"42",X"02",X"02",X"02",X"37",X"38",X"42",X"C1",X"44",X"05",X"81",X"02",X"01",
		X"02",X"02",X"02",X"3F",X"3E",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"02",X"37",X"38",
		X"04",X"42",X"C1",X"44",X"05",X"81",X"02",X"00",X"02",X"02",X"3F",X"3E",X"33",X"42",X"C1",X"44",
		X"05",X"81",X"42",X"02",X"02",X"37",X"38",X"04",X"30",X"02",X"C1",X"44",X"05",X"81",X"02",X"02",
		X"02",X"3F",X"3E",X"33",X"34",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",X"37",X"38",X"04",X"30",
		X"31",X"02",X"C1",X"44",X"05",X"81",X"02",X"02",X"3F",X"3E",X"33",X"34",X"02",X"02",X"C1",X"44",
		X"05",X"81",X"01",X"37",X"38",X"04",X"30",X"31",X"02",X"42",X"C1",X"44",X"05",X"81",X"02",X"3F",
		X"3E",X"33",X"34",X"02",X"02",X"42",X"C1",X"44",X"05",X"81",X"37",X"38",X"04",X"30",X"31",X"40",
		X"02",X"42",X"C1",X"44",X"05",X"81",X"3F",X"3E",X"33",X"34",X"02",X"42",X"42",X"42",X"C1",X"44",
		X"05",X"78",X"38",X"04",X"30",X"31",X"02",X"ED",X"AD",X"02",X"C1",X"44",X"07",X"33",X"34",X"02",
		X"02",X"02",X"02",X"42",X"C1",X"44",X"07",X"30",X"31",X"42",X"02",X"02",X"41",X"02",X"C1",X"44",
		X"06",X"33",X"34",X"02",X"ED",X"AD",X"02",X"02",X"02",X"C1",X"44",X"06",X"30",X"31",X"42",X"42",
		X"02",X"01",X"02",X"42",X"C1",X"44",X"05",X"33",X"34",X"02",X"01",X"02",X"02",X"02",X"02",X"42",
		X"C1",X"44",X"05",X"30",X"31",X"02",X"42",X"02",X"ED",X"AD",X"02",X"42",X"C1",X"44",X"05",X"81",
		X"42",X"ED",X"AD",X"02",X"02",X"42",X"42",X"42",X"C1",X"44",X"05",X"81",X"02",X"02",X"02",X"42",
		X"02",X"ED",X"AD",X"02",X"C1",X"44",X"05",X"81",X"02",X"40",X"02",X"02",X"02",X"02",X"02",X"42",
		X"C1",X"44",X"05",X"81",X"02",X"02",X"ED",X"AD",X"02",X"02",X"02",X"02",X"C1",X"44",X"05",X"81",
		X"02",X"02",X"02",X"42",X"42",X"01",X"02",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"0C",X"0C",X"71",X"21",X"6D",X"F3",X"35",X"C2",X"B6",X"9D",X"3A",X"2F",X"F0",X"3D",X"32",X"2F",
		X"F0",X"FE",X"01",X"28",X"20",X"38",X"33",X"21",X"98",X"E8",X"11",X"F8",X"9C",X"CD",X"18",X"3F",
		X"21",X"D8",X"E8",X"11",X"0D",X"9D",X"CD",X"18",X"3F",X"21",X"18",X"E9",X"11",X"22",X"9D",X"CD",
		X"18",X"3F",X"C3",X"B6",X"9D",X"21",X"98",X"E8",X"CD",X"15",X"3F",X"21",X"D8",X"E8",X"CD",X"15",
		X"3F",X"21",X"18",X"E9",X"CD",X"15",X"3F",X"C3",X"B6",X"9D",X"CD",X"BC",X"89",X"CD",X"3A",X"3D",
		X"C9",X"21",X"82",X"F3",X"11",X"76",X"F3",X"7E",X"12",X"13",X"23",X"06",X"03",X"7E",X"CB",X"27",
		X"CB",X"27",X"CB",X"27",X"CB",X"27",X"23",X"B6",X"12",X"13",X"23",X"10",X"F0",X"C9",X"DD",X"21",
		X"5B",X"F4",X"21",X"60",X"F3",X"3E",X"0A",X"96",X"28",X"1A",X"47",X"11",X"FD",X"FF",X"DD",X"19",
		X"DD",X"7E",X"00",X"DD",X"77",X"03",X"DD",X"7E",X"01",X"DD",X"77",X"04",X"DD",X"7E",X"02",X"DD",
		X"77",X"05",X"10",X"EA",X"FD",X"21",X"90",X"E9",X"06",X"03",X"FD",X"7E",X"00",X"B7",X"20",X"02",
		X"3E",X"20",X"DD",X"77",X"00",X"DD",X"23",X"FD",X"2B",X"FD",X"2B",X"10",X"ED",X"C9",X"11",X"63",
		X"A1",X"21",X"75",X"E9",X"CD",X"18",X"3F",X"11",X"70",X"A1",X"21",X"D5",X"E9",X"CD",X"18",X"3F",
		X"CD",X"51",X"A0",X"0E",X"65",X"DD",X"21",X"F6",X"F5",X"21",X"76",X"F3",X"06",X"04",X"DD",X"E5",
		X"7E",X"DD",X"BE",X"00",X"38",X"2B",X"20",X"05",X"23",X"DD",X"23",X"10",X"F3",X"DD",X"E1",X"79",
		X"FE",X"65",X"28",X"10",X"DD",X"E5",X"06",X"04",X"DD",X"7E",X"00",X"DD",X"77",X"04",X"DD",X"23",
		X"10",X"F6",X"DD",X"E1",X"11",X"FC",X"FF",X"DD",X"19",X"0D",X"79",X"FE",X"01",X"20",X"CA",X"18",
		X"1D",X"DD",X"E1",X"79",X"FE",X"65",X"38",X"16",X"32",X"60",X"F3",X"11",X"7D",X"A1",X"21",X"35",
		X"EA",X"CD",X"18",X"3F",X"11",X"8C",X"A1",X"21",X"95",X"EA",X"CD",X"18",X"3F",X"C9",X"32",X"60",
		X"F3",X"21",X"76",X"F3",X"06",X"04",X"7E",X"DD",X"77",X"04",X"23",X"DD",X"23",X"10",X"F7",X"21",
		X"64",X"F3",X"36",X"20",X"06",X"20",X"3A",X"60",X"F3",X"FE",X"64",X"38",X"06",X"36",X"31",X"D6",
		X"64",X"06",X"30",X"23",X"FE",X"0A",X"38",X"09",X"06",X"30",X"D6",X"0A",X"04",X"FE",X"0A",X"30",
		X"F9",X"70",X"23",X"C6",X"30",X"77",X"23",X"36",X"00",X"11",X"64",X"F3",X"21",X"30",X"EA",X"CD",
		X"18",X"3F",X"C9",X"20",X"20",X"59",X"4F",X"55",X"52",X"20",X"53",X"43",X"4F",X"52",X"45",X"00",
		X"20",X"20",X"52",X"41",X"4E",X"4B",X"49",X"4E",X"47",X"20",X"49",X"53",X"00",X"4E",X"4F",X"54",
		X"20",X"49",X"4E",X"20",X"54",X"48",X"45",X"20",X"54",X"4F",X"50",X"00",X"20",X"20",X"31",X"30",
		X"30",X"20",X"53",X"43",X"4F",X"52",X"45",X"53",X"00",X"21",X"0E",X"F6",X"DD",X"21",X"27",X"A2",
		X"06",X"09",X"3A",X"8B",X"F3",X"DD",X"BE",X"00",X"38",X"14",X"20",X"0A",X"3A",X"8C",X"F3",X"DD",
		X"BE",X"01",X"38",X"0A",X"28",X"08",X"23",X"23",X"DD",X"23",X"DD",X"23",X"10",X"E4",X"34",X"20",
		X"2B",X"23",X"34",X"20",X"27",X"35",X"2B",X"35",X"06",X"0A",X"11",X"00",X"FF",X"DD",X"21",X"0E",
		X"F6",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"7C",X"B7",X"28",X"03",X"19",X"18",X"02",X"2E",X"00",
		X"DD",X"75",X"00",X"DD",X"74",X"01",X"DD",X"23",X"DD",X"23",X"10",X"E5",X"21",X"5E",X"F4",X"3A",
		X"8B",X"F3",X"BE",X"38",X"15",X"20",X"07",X"23",X"3A",X"8C",X"F3",X"BE",X"38",X"0C",X"3A",X"8B",
		X"F3",X"32",X"5E",X"F4",X"3A",X"8C",X"F3",X"32",X"5F",X"F4",X"21",X"60",X"F4",X"3A",X"8B",X"F3",
		X"BE",X"38",X"07",X"C0",X"3A",X"8C",X"F3",X"23",X"BE",X"D0",X"3A",X"8B",X"F3",X"32",X"60",X"F4",
		X"3A",X"8C",X"F3",X"32",X"61",X"F4",X"C9",X"01",X"30",X"02",X"00",X"02",X"30",X"03",X"00",X"04",
		X"00",X"05",X"00",X"07",X"00",X"10",X"00",X"15",X"00",X"21",X"FA",X"F5",X"DD",X"21",X"F0",X"A2",
		X"06",X"09",X"3A",X"77",X"F3",X"DD",X"BE",X"00",X"38",X"20",X"20",X"14",X"3A",X"78",X"F3",X"DD",
		X"BE",X"01",X"38",X"16",X"20",X"0A",X"3A",X"79",X"F3",X"DD",X"BE",X"02",X"38",X"0C",X"28",X"0A",
		X"23",X"23",X"DD",X"23",X"DD",X"23",X"DD",X"23",X"10",X"D8",X"34",X"20",X"2B",X"23",X"34",X"20",
		X"27",X"35",X"2B",X"35",X"06",X"0A",X"11",X"00",X"FF",X"DD",X"21",X"0E",X"F6",X"DD",X"6E",X"00",
		X"DD",X"66",X"01",X"7C",X"B7",X"28",X"03",X"19",X"18",X"02",X"2E",X"00",X"DD",X"75",X"00",X"DD",
		X"74",X"01",X"DD",X"23",X"DD",X"23",X"10",X"E5",X"21",X"62",X"F4",X"3A",X"77",X"F3",X"BE",X"38",
		X"24",X"20",X"10",X"23",X"3A",X"78",X"F3",X"BE",X"38",X"1B",X"20",X"07",X"23",X"3A",X"79",X"F3",
		X"BE",X"38",X"12",X"3A",X"77",X"F3",X"32",X"62",X"F4",X"3A",X"78",X"F3",X"32",X"63",X"F4",X"3A",
		X"79",X"F3",X"32",X"64",X"F4",X"21",X"66",X"F4",X"3A",X"77",X"F3",X"BE",X"38",X"0F",X"C0",X"3A",
		X"78",X"F3",X"23",X"BE",X"38",X"07",X"C0",X"23",X"3A",X"79",X"F3",X"BE",X"D0",X"3A",X"77",X"F3",
		X"32",X"66",X"F4",X"3A",X"78",X"F3",X"32",X"67",X"F4",X"3A",X"79",X"F3",X"32",X"68",X"F4",X"C9",
		X"00",X"50",X"00",X"01",X"00",X"00",X"01",X"32",X"00",X"02",X"00",X"00",X"02",X"50",X"00",X"03",
		X"00",X"00",X"05",X"00",X"00",X"07",X"50",X"00",X"10",X"00",X"00",X"CD",X"25",X"3D",X"21",X"A6",
		X"F0",X"36",X"13",X"3E",X"78",X"32",X"1A",X"F4",X"21",X"00",X"F8",X"36",X"FE",X"0E",X"02",X"CD",
		X"4E",X"3D",X"21",X"2D",X"A4",X"22",X"00",X"F1",X"3E",X"08",X"32",X"02",X"F1",X"3E",X"01",X"32",
		X"16",X"F4",X"AF",X"32",X"01",X"F4",X"DB",X"01",X"2F",X"E6",X"04",X"32",X"04",X"F1",X"CD",X"3A",
		X"3D",X"0E",X"02",X"CD",X"4E",X"3D",X"CD",X"67",X"09",X"CD",X"4C",X"09",X"CD",X"C3",X"A3",X"DD",
		X"2A",X"00",X"F1",X"DD",X"7E",X"07",X"32",X"06",X"F8",X"CD",X"EC",X"A3",X"DB",X"00",X"2F",X"E6",
		X"80",X"CA",X"00",X"00",X"CD",X"F9",X"3C",X"CD",X"77",X"A3",X"CD",X"EC",X"A3",X"CD",X"AB",X"A3",
		X"28",X"EA",X"CD",X"11",X"A4",X"18",X"94",X"21",X"02",X"F1",X"35",X"C0",X"36",X"08",X"21",X"03",
		X"F1",X"DD",X"2A",X"00",X"F1",X"DB",X"01",X"2F",X"E6",X"08",X"28",X"0C",X"7E",X"B7",X"28",X"03",
		X"35",X"18",X"05",X"DD",X"7E",X"06",X"3D",X"77",X"DB",X"01",X"2F",X"E6",X"01",X"C8",X"DD",X"46",
		X"06",X"05",X"7E",X"B8",X"30",X"02",X"34",X"C9",X"36",X"00",X"C9",X"3A",X"04",X"F1",X"47",X"DB",
		X"01",X"2F",X"E6",X"04",X"32",X"04",X"F1",X"B7",X"28",X"04",X"78",X"B7",X"28",X"02",X"AF",X"C9",
		X"F6",X"01",X"C9",X"DD",X"2A",X"00",X"F1",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E5",X"DD",X"E1",
		X"DD",X"6E",X"00",X"DD",X"66",X"01",X"7C",X"B5",X"C8",X"DD",X"5E",X"02",X"DD",X"56",X"03",X"CD",
		X"18",X"3F",X"11",X"04",X"00",X"DD",X"19",X"CD",X"F9",X"3C",X"18",X"E4",X"DD",X"2A",X"00",X"F1",
		X"DD",X"6E",X"02",X"DD",X"66",X"03",X"16",X"00",X"3A",X"03",X"F1",X"5F",X"19",X"19",X"DD",X"21",
		X"04",X"F8",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"03",X"3E",X"34",X"DD",X"77",X"02",
		X"C9",X"DD",X"2A",X"00",X"F1",X"DD",X"6E",X"04",X"DD",X"66",X"05",X"16",X"00",X"3A",X"03",X"F1",
		X"5F",X"19",X"19",X"E5",X"DD",X"E1",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E9",X"59",X"A4",X"35",
		X"A4",X"47",X"A4",X"09",X"34",X"30",X"24",X"30",X"34",X"30",X"44",X"30",X"54",X"30",X"64",X"30",
		X"74",X"30",X"84",X"30",X"94",X"30",X"A4",X"16",X"08",X"92",X"A5",X"A3",X"B2",X"10",X"A9",X"FA",
		X"B5",X"E7",X"AD",X"95",X"13",X"70",X"0B",X"DC",X"AE",X"79",X"E8",X"93",X"A4",X"B7",X"E8",X"A7",
		X"A4",X"F7",X"E8",X"BA",X"A4",X"37",X"E9",X"C3",X"A4",X"77",X"E9",X"D2",X"A4",X"B7",X"E9",X"E0",
		X"A4",X"F7",X"E9",X"F0",X"A4",X"37",X"EA",X"FF",X"A4",X"77",X"EA",X"08",X"A5",X"B7",X"EA",X"17",
		X"A5",X"1B",X"EB",X"29",X"A5",X"3B",X"EB",X"43",X"A5",X"7B",X"EB",X"5F",X"A5",X"9B",X"EB",X"7A",
		X"A5",X"00",X"00",X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"44",X"45",X"53",X"49",X"52",X"45",
		X"44",X"20",X"54",X"45",X"53",X"54",X"00",X"31",X"20",X"53",X"45",X"4C",X"46",X"20",X"44",X"49",
		X"41",X"47",X"4E",X"4F",X"53",X"54",X"49",X"43",X"53",X"00",X"32",X"20",X"53",X"4F",X"55",X"4E",
		X"44",X"53",X"00",X"33",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"49",X"4E",X"50",X"55",
		X"54",X"00",X"34",X"20",X"42",X"4F",X"4F",X"4B",X"4B",X"45",X"45",X"50",X"49",X"4E",X"47",X"00",
		X"35",X"20",X"4D",X"41",X"43",X"48",X"49",X"4E",X"45",X"20",X"53",X"45",X"54",X"55",X"50",X"00",
		X"36",X"20",X"43",X"48",X"41",X"4E",X"4E",X"45",X"4C",X"20",X"54",X"45",X"53",X"54",X"00",X"37",
		X"20",X"50",X"52",X"45",X"53",X"45",X"54",X"00",X"38",X"20",X"47",X"52",X"49",X"44",X"20",X"44",
		X"49",X"53",X"50",X"4C",X"41",X"59",X"00",X"39",X"20",X"50",X"4F",X"54",X"20",X"43",X"41",X"4C",
		X"49",X"42",X"52",X"41",X"54",X"49",X"4F",X"4E",X"00",X"50",X"4F",X"53",X"49",X"54",X"49",X"4F",
		X"4E",X"20",X"43",X"55",X"52",X"53",X"4F",X"52",X"20",X"55",X"53",X"49",X"4E",X"47",X"20",X"54",
		X"48",X"45",X"00",X"53",X"4D",X"4F",X"4B",X"45",X"20",X"41",X"4E",X"44",X"20",X"4F",X"49",X"4C",
		X"20",X"54",X"48",X"55",X"4D",X"42",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"53",X"00",X"55",
		X"53",X"45",X"20",X"54",X"48",X"45",X"20",X"57",X"45",X"41",X"50",X"4F",X"4E",X"53",X"20",X"56",
		X"41",X"4E",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"54",X"4F",X"20",X"53",X"45",X"4C",
		X"45",X"43",X"54",X"20",X"41",X"20",X"54",X"45",X"53",X"54",X"20",X"4F",X"50",X"54",X"49",X"4F",
		X"4E",X"00",X"21",X"A6",X"F0",X"36",X"11",X"21",X"60",X"A6",X"22",X"00",X"F1",X"21",X"C8",X"A8",
		X"22",X"07",X"F1",X"3E",X"08",X"AF",X"32",X"03",X"F1",X"32",X"05",X"F1",X"CD",X"67",X"09",X"CD",
		X"4C",X"09",X"CD",X"3A",X"3D",X"CD",X"F9",X"3C",X"CD",X"85",X"0B",X"0E",X"02",X"CD",X"4E",X"3D",
		X"CD",X"F9",X"3C",X"0E",X"02",X"CD",X"4E",X"3D",X"CD",X"C3",X"A3",X"DD",X"2A",X"00",X"F1",X"DD",
		X"7E",X"07",X"32",X"06",X"F8",X"3A",X"05",X"F1",X"B7",X"20",X"1D",X"DB",X"00",X"2F",X"E6",X"80",
		X"28",X"16",X"CD",X"F9",X"3C",X"CD",X"77",X"A3",X"CD",X"EC",X"A3",X"CD",X"AB",X"A3",X"28",X"E5",
		X"CD",X"F8",X"A5",X"CD",X"11",X"A4",X"18",X"DD",X"21",X"A6",X"F0",X"36",X"13",X"C9",X"2A",X"07",
		X"F1",X"16",X"00",X"3A",X"03",X"F1",X"D6",X"02",X"5F",X"19",X"19",X"19",X"E5",X"DD",X"E1",X"DD",
		X"4E",X"00",X"CD",X"4E",X"3D",X"DD",X"46",X"01",X"04",X"CD",X"F9",X"3C",X"10",X"FB",X"DD",X"7E",
		X"02",X"B7",X"FA",X"28",X"A6",X"20",X"05",X"C9",X"0E",X"02",X"18",X"01",X"4F",X"CD",X"4E",X"3D",
		X"C9",X"3E",X"02",X"32",X"03",X"F1",X"3A",X"03",X"F1",X"DD",X"2A",X"00",X"F1",X"DD",X"BE",X"06",
		X"30",X"13",X"CD",X"EC",X"A3",X"06",X"0A",X"CD",X"F9",X"3C",X"10",X"FB",X"CD",X"FE",X"A5",X"21",
		X"03",X"F1",X"34",X"18",X"E1",X"AF",X"32",X"03",X"F1",X"C9",X"3E",X"01",X"32",X"05",X"F1",X"C9",
		X"9C",X"A6",X"68",X"A6",X"94",X"A8",X"1A",X"34",X"28",X"1C",X"28",X"24",X"28",X"2C",X"28",X"34",
		X"28",X"3C",X"28",X"44",X"28",X"4C",X"28",X"54",X"28",X"5C",X"28",X"64",X"28",X"6C",X"28",X"74",
		X"28",X"7C",X"28",X"84",X"28",X"8C",X"28",X"94",X"28",X"9C",X"28",X"A4",X"28",X"AC",X"28",X"B4",
		X"28",X"BC",X"28",X"C4",X"28",X"CC",X"28",X"D4",X"28",X"DC",X"28",X"E4",X"57",X"E8",X"0A",X"A7",
		X"97",X"E8",X"19",X"A7",X"B7",X"E8",X"26",X"A7",X"D7",X"E8",X"2D",X"A7",X"F7",X"E8",X"34",X"A7",
		X"17",X"E9",X"41",X"A7",X"37",X"E9",X"48",X"A7",X"57",X"E9",X"54",X"A7",X"77",X"E9",X"61",X"A7",
		X"97",X"E9",X"6D",X"A7",X"B8",X"E9",X"7C",X"A7",X"D8",X"E9",X"8C",X"A7",X"F8",X"E9",X"9E",X"A7",
		X"18",X"EA",X"AE",X"A7",X"38",X"EA",X"BB",X"A7",X"58",X"EA",X"CB",X"A7",X"78",X"EA",X"D9",X"A7",
		X"98",X"EA",X"E9",X"A7",X"B8",X"EA",X"FF",X"A7",X"D8",X"EA",X"0E",X"A8",X"F8",X"EA",X"25",X"A8",
		X"18",X"EB",X"39",X"A8",X"38",X"EB",X"45",X"A8",X"58",X"EB",X"57",X"A8",X"78",X"EB",X"66",X"A8",
		X"98",X"EB",X"76",X"A8",X"B8",X"EB",X"89",X"A8",X"00",X"00",X"53",X"45",X"4C",X"45",X"43",X"54",
		X"20",X"41",X"20",X"53",X"4F",X"55",X"4E",X"44",X"00",X"31",X"20",X"41",X"4C",X"4C",X"20",X"53",
		X"4F",X"55",X"4E",X"44",X"53",X"00",X"32",X"20",X"45",X"58",X"49",X"54",X"00",X"33",X"20",X"43",
		X"4F",X"49",X"4E",X"00",X"34",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"42",X"41",X"53",X"45",
		X"00",X"35",X"20",X"54",X"49",X"4C",X"54",X"00",X"36",X"20",X"42",X"4F",X"4D",X"42",X"20",X"46",
		X"41",X"4C",X"4C",X"00",X"37",X"20",X"45",X"58",X"50",X"4C",X"4F",X"53",X"49",X"4F",X"4E",X"20",
		X"00",X"38",X"20",X"43",X"41",X"52",X"20",X"43",X"52",X"41",X"53",X"48",X"00",X"39",X"20",X"53",
		X"48",X"4F",X"54",X"47",X"55",X"4E",X"20",X"46",X"49",X"52",X"45",X"00",X"31",X"30",X"20",X"43",
		X"41",X"52",X"20",X"4F",X"46",X"46",X"20",X"52",X"4F",X"41",X"44",X"00",X"31",X"31",X"20",X"53",
		X"54",X"41",X"4C",X"4C",X"45",X"44",X"20",X"45",X"4E",X"47",X"49",X"4E",X"45",X"00",X"31",X"32",
		X"20",X"4D",X"41",X"43",X"48",X"49",X"4E",X"45",X"20",X"47",X"55",X"4E",X"53",X"00",X"31",X"33",
		X"20",X"4F",X"49",X"4C",X"20",X"53",X"4C",X"49",X"43",X"4B",X"00",X"31",X"34",X"20",X"53",X"4D",
		X"4F",X"4B",X"45",X"20",X"53",X"43",X"52",X"45",X"45",X"4E",X"00",X"31",X"35",X"20",X"54",X"49",
		X"52",X"45",X"20",X"43",X"48",X"49",X"52",X"50",X"00",X"31",X"36",X"20",X"54",X"49",X"52",X"45",
		X"20",X"53",X"4C",X"41",X"53",X"48",X"45",X"52",X"00",X"31",X"37",X"20",X"48",X"45",X"4C",X"49",
		X"43",X"4F",X"50",X"54",X"45",X"52",X"20",X"46",X"41",X"44",X"45",X"20",X"49",X"4E",X"00",X"31",
		X"38",X"20",X"48",X"45",X"4C",X"49",X"43",X"4F",X"50",X"54",X"45",X"52",X"20",X"00",X"31",X"39",
		X"20",X"48",X"45",X"4C",X"49",X"43",X"4F",X"50",X"54",X"45",X"52",X"20",X"46",X"41",X"44",X"45",
		X"20",X"4F",X"55",X"54",X"00",X"32",X"30",X"20",X"48",X"45",X"4C",X"49",X"43",X"4F",X"50",X"54",
		X"45",X"52",X"20",X"43",X"52",X"41",X"53",X"48",X"00",X"32",X"31",X"20",X"54",X"55",X"47",X"20",
		X"42",X"4F",X"41",X"54",X"00",X"32",X"32",X"20",X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"20",
		X"4C",X"41",X"55",X"4E",X"43",X"48",X"00",X"32",X"33",X"20",X"43",X"41",X"52",X"20",X"53",X"50",
		X"4C",X"41",X"53",X"48",X"20",X"00",X"32",X"34",X"20",X"43",X"41",X"52",X"20",X"53",X"50",X"49",
		X"4E",X"20",X"4F",X"55",X"54",X"00",X"32",X"35",X"20",X"42",X"55",X"4C",X"4C",X"45",X"54",X"20",
		X"52",X"49",X"43",X"4F",X"43",X"48",X"45",X"54",X"00",X"32",X"36",X"20",X"54",X"4F",X"52",X"50",
		X"45",X"44",X"4F",X"00",X"31",X"A6",X"5A",X"A6",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",
		X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",
		X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",
		X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"FE",X"A5",X"0C",X"1E",X"FF",X"0B",X"1E",X"00",X"09",X"3C",
		X"FF",X"0D",X"50",X"00",X"19",X"3C",X"1A",X"13",X"28",X"14",X"1B",X"1E",X"1C",X"1D",X"1E",X"00",
		X"1F",X"28",X"20",X"22",X"28",X"23",X"24",X"3C",X"21",X"25",X"B0",X"00",X"26",X"28",X"00",X"27",
		X"28",X"28",X"29",X"3C",X"2A",X"2B",X"3C",X"2A",X"2C",X"3C",X"2A",X"15",X"3C",X"16",X"4F",X"3C",
		X"00",X"30",X"28",X"00",X"33",X"28",X"00",X"35",X"28",X"00",X"37",X"28",X"00",X"2F",X"50",X"4C",
		X"21",X"5B",X"A9",X"22",X"00",X"F1",X"3E",X"08",X"AF",X"32",X"03",X"F1",X"32",X"05",X"F1",X"CD",
		X"67",X"09",X"CD",X"4C",X"09",X"CD",X"3A",X"3D",X"0E",X"02",X"CD",X"4E",X"3D",X"CD",X"C3",X"A3",
		X"DD",X"2A",X"00",X"F1",X"DD",X"7E",X"07",X"32",X"06",X"F8",X"CD",X"3A",X"AA",X"3A",X"05",X"F1",
		X"B7",X"C0",X"DB",X"00",X"2F",X"E6",X"80",X"C8",X"CD",X"F9",X"3C",X"CD",X"77",X"A3",X"CD",X"EC",
		X"A3",X"CD",X"AB",X"A3",X"28",X"E7",X"CD",X"11",X"A4",X"18",X"C4",X"69",X"A9",X"63",X"A9",X"34",
		X"AA",X"03",X"34",X"98",X"86",X"98",X"96",X"98",X"A6",X"7C",X"E8",X"A3",X"A9",X"BB",X"E8",X"BB",
		X"A9",X"FB",X"E8",X"CA",X"A9",X"3B",X"E9",X"D9",X"A9",X"7B",X"E9",X"E6",X"A9",X"BB",X"E9",X"F4",
		X"A9",X"FB",X"E9",X"02",X"AA",X"3B",X"EA",X"16",X"AA",X"7B",X"EA",X"22",X"AA",X"BB",X"EA",X"2F",
		X"AA",X"FB",X"EA",X"29",X"A5",X"1B",X"EB",X"43",X"A5",X"5B",X"EB",X"5F",X"A5",X"7B",X"EB",X"7A",
		X"A5",X"00",X"00",X"53",X"45",X"4C",X"45",X"43",X"54",X"20",X"41",X"20",X"52",X"45",X"50",X"4F",
		X"52",X"54",X"20",X"4F",X"52",X"20",X"45",X"58",X"49",X"54",X"00",X"43",X"48",X"55",X"54",X"45",
		X"20",X"20",X"31",X"20",X"43",X"4F",X"49",X"4E",X"53",X"00",X"43",X"48",X"55",X"54",X"45",X"20",
		X"20",X"32",X"20",X"43",X"4F",X"49",X"4E",X"53",X"00",X"4C",X"4F",X"4E",X"47",X"45",X"53",X"54",
		X"20",X"47",X"41",X"4D",X"45",X"00",X"53",X"48",X"4F",X"52",X"54",X"45",X"53",X"54",X"20",X"47",
		X"41",X"4D",X"45",X"00",X"48",X"49",X"47",X"48",X"45",X"53",X"54",X"20",X"53",X"43",X"4F",X"52",
		X"45",X"00",X"4C",X"4F",X"57",X"45",X"53",X"54",X"20",X"53",X"43",X"4F",X"52",X"45",X"00",X"42",
		X"55",X"59",X"20",X"49",X"4E",X"00",X"54",X"49",X"4D",X"45",X"20",X"52",X"45",X"50",X"4F",X"52",
		X"54",X"00",X"53",X"43",X"4F",X"52",X"45",X"20",X"52",X"45",X"50",X"4F",X"52",X"54",X"00",X"45",
		X"58",X"49",X"54",X"00",X"26",X"AB",X"92",X"AC",X"5A",X"A6",X"2A",X"22",X"F6",X"DD",X"21",X"19",
		X"F1",X"CD",X"CA",X"AA",X"06",X"05",X"0E",X"00",X"1E",X"01",X"DD",X"21",X"AA",X"E8",X"21",X"19",
		X"F1",X"CD",X"DA",X"AA",X"2A",X"24",X"F6",X"DD",X"21",X"19",X"F1",X"CD",X"CA",X"AA",X"06",X"05",
		X"0E",X"00",X"1E",X"01",X"DD",X"21",X"EA",X"E8",X"21",X"19",X"F1",X"CD",X"DA",X"AA",X"21",X"5E",
		X"F4",X"DD",X"21",X"2A",X"E9",X"CD",X"10",X"AB",X"21",X"60",X"F4",X"DD",X"21",X"6A",X"E9",X"CD",
		X"10",X"AB",X"06",X"06",X"0E",X"00",X"DD",X"21",X"AB",X"E9",X"21",X"62",X"F4",X"CD",X"D8",X"AA",
		X"06",X"06",X"0E",X"00",X"DD",X"21",X"EB",X"E9",X"21",X"66",X"F4",X"C3",X"D8",X"AA",X"06",X"03",
		X"AF",X"DD",X"77",X"00",X"DD",X"77",X"01",X"DD",X"77",X"02",X"FD",X"5E",X"00",X"FD",X"23",X"FD",
		X"56",X"00",X"FD",X"23",X"B7",X"ED",X"52",X"38",X"0B",X"DD",X"7E",X"00",X"C6",X"01",X"27",X"DD",
		X"77",X"00",X"18",X"F0",X"19",X"DD",X"23",X"10",X"E1",X"C9",X"FD",X"21",X"D2",X"AA",X"CD",X"9E",
		X"AA",X"C9",X"10",X"27",X"64",X"00",X"01",X"00",X"1E",X"00",X"7B",X"B7",X"7E",X"28",X"05",X"1E",
		X"00",X"23",X"18",X"06",X"1F",X"1F",X"1F",X"1F",X"1E",X"01",X"E6",X"0F",X"05",X"20",X"02",X"0E",
		X"01",X"04",X"C6",X"30",X"FE",X"30",X"20",X"0A",X"0C",X"0D",X"20",X"07",X"DD",X"36",X"00",X"00",
		X"18",X"04",X"4F",X"DD",X"77",X"00",X"D5",X"11",X"FF",X"FF",X"DD",X"19",X"D1",X"10",X"CB",X"C9",
		X"01",X"02",X"02",X"CD",X"D8",X"AA",X"DD",X"36",X"00",X"00",X"01",X"FF",X"FF",X"DD",X"09",X"01",
		X"02",X"02",X"CD",X"D8",X"AA",X"C9",X"CD",X"67",X"09",X"CD",X"4C",X"09",X"CD",X"3A",X"3D",X"DD",
		X"21",X"7C",X"AB",X"CD",X"D0",X"A3",X"06",X"0A",X"21",X"0E",X"F6",X"FD",X"21",X"7E",X"AC",X"5E",
		X"23",X"56",X"23",X"E5",X"C5",X"FD",X"E5",X"EB",X"DD",X"21",X"19",X"F1",X"CD",X"CA",X"AA",X"06",
		X"05",X"0E",X"00",X"1E",X"01",X"21",X"19",X"F1",X"FD",X"E1",X"FD",X"5E",X"00",X"FD",X"56",X"01",
		X"D5",X"DD",X"E1",X"FD",X"23",X"FD",X"23",X"CD",X"DA",X"AA",X"C1",X"E1",X"10",X"D1",X"CD",X"F9",
		X"3C",X"CD",X"AB",X"A3",X"C0",X"DB",X"00",X"E6",X"80",X"C0",X"18",X"F2",X"75",X"E8",X"B2",X"AB",
		X"BB",X"E8",X"BE",X"AB",X"FB",X"E8",X"CD",X"AB",X"3B",X"E9",X"DC",X"AB",X"7B",X"E9",X"EB",X"AB",
		X"BB",X"E9",X"FA",X"AB",X"FB",X"E9",X"09",X"AC",X"3B",X"EA",X"18",X"AC",X"7B",X"EA",X"27",X"AC",
		X"BB",X"EA",X"36",X"AC",X"FB",X"EA",X"45",X"AC",X"5B",X"EB",X"54",X"AC",X"9B",X"EB",X"6A",X"AC",
		X"00",X"00",X"54",X"49",X"4D",X"45",X"20",X"52",X"45",X"50",X"4F",X"52",X"54",X"00",X"20",X"20",
		X"30",X"20",X"54",X"4F",X"20",X"20",X"39",X"30",X"20",X"53",X"45",X"43",X"00",X"20",X"39",X"30",
		X"20",X"54",X"4F",X"20",X"31",X"32",X"30",X"20",X"53",X"45",X"43",X"00",X"31",X"32",X"30",X"20",
		X"54",X"4F",X"20",X"31",X"35",X"30",X"20",X"53",X"45",X"43",X"00",X"31",X"35",X"30",X"20",X"54",
		X"4F",X"20",X"31",X"38",X"30",X"20",X"53",X"45",X"43",X"00",X"20",X"20",X"33",X"20",X"54",X"4F",
		X"20",X"20",X"20",X"34",X"20",X"4D",X"49",X"4E",X"00",X"20",X"20",X"34",X"20",X"54",X"4F",X"20",
		X"20",X"20",X"35",X"20",X"4D",X"49",X"4E",X"00",X"20",X"20",X"35",X"20",X"54",X"4F",X"20",X"20",
		X"20",X"37",X"20",X"4D",X"49",X"4E",X"00",X"20",X"20",X"37",X"20",X"54",X"4F",X"20",X"20",X"31",
		X"30",X"20",X"4D",X"49",X"4E",X"00",X"20",X"31",X"30",X"20",X"54",X"4F",X"20",X"20",X"31",X"35",
		X"20",X"4D",X"49",X"4E",X"00",X"20",X"20",X"20",X"4F",X"56",X"45",X"52",X"20",X"31",X"35",X"20",
		X"4D",X"49",X"4E",X"00",X"50",X"52",X"45",X"53",X"53",X"20",X"54",X"48",X"45",X"20",X"57",X"45",
		X"41",X"50",X"4F",X"4E",X"53",X"20",X"56",X"41",X"4E",X"00",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"20",X"54",X"4F",X"20",X"45",X"58",X"49",X"54",X"20",X"54",X"45",X"53",X"54",X"00",X"A9",X"E8",
		X"E9",X"E8",X"29",X"E9",X"69",X"E9",X"A9",X"E9",X"E9",X"E9",X"29",X"EA",X"69",X"EA",X"A9",X"EA",
		X"E9",X"EA",X"CD",X"67",X"09",X"CD",X"4C",X"09",X"CD",X"3A",X"3D",X"DD",X"21",X"E6",X"AC",X"CD",
		X"D0",X"A3",X"06",X"0A",X"21",X"FA",X"F5",X"FD",X"21",X"D3",X"AD",X"5E",X"23",X"56",X"23",X"E5",
		X"C5",X"FD",X"E5",X"EB",X"DD",X"21",X"19",X"F1",X"CD",X"CA",X"AA",X"06",X"06",X"0E",X"00",X"21",
		X"19",X"F1",X"FD",X"E1",X"FD",X"5E",X"00",X"FD",X"56",X"01",X"D5",X"DD",X"E1",X"FD",X"23",X"FD",
		X"23",X"CD",X"D8",X"AA",X"C1",X"E1",X"10",X"D3",X"CD",X"F9",X"3C",X"CD",X"AB",X"A3",X"C0",X"DB",
		X"00",X"E6",X"80",X"C0",X"18",X"F2",X"55",X"E8",X"1C",X"AD",X"BB",X"E8",X"29",X"AD",X"FB",X"E8",
		X"3A",X"AD",X"3B",X"E9",X"4B",X"AD",X"7B",X"E9",X"5C",X"AD",X"BB",X"E9",X"6D",X"AD",X"FB",X"E9",
		X"7E",X"AD",X"3B",X"EA",X"8F",X"AD",X"7B",X"EA",X"A0",X"AD",X"BB",X"EA",X"B1",X"AD",X"FB",X"EA",
		X"C2",X"AD",X"5B",X"EB",X"54",X"AC",X"9B",X"EB",X"6A",X"AC",X"00",X"00",X"53",X"43",X"4F",X"52",
		X"45",X"20",X"52",X"45",X"50",X"4F",X"52",X"54",X"00",X"20",X"20",X"20",X"20",X"20",X"30",X"20",
		X"54",X"4F",X"20",X"20",X"20",X"35",X"30",X"30",X"30",X"00",X"20",X"20",X"35",X"30",X"30",X"30",
		X"20",X"54",X"4F",X"20",X"20",X"31",X"30",X"30",X"30",X"30",X"00",X"20",X"31",X"30",X"30",X"30",
		X"30",X"20",X"54",X"4F",X"20",X"20",X"31",X"35",X"30",X"30",X"30",X"00",X"20",X"31",X"35",X"30",
		X"30",X"30",X"20",X"54",X"4F",X"20",X"20",X"32",X"30",X"30",X"30",X"30",X"00",X"20",X"32",X"30",
		X"30",X"30",X"30",X"20",X"54",X"4F",X"20",X"20",X"32",X"35",X"30",X"30",X"30",X"00",X"20",X"32",
		X"35",X"30",X"30",X"30",X"20",X"54",X"4F",X"20",X"20",X"33",X"30",X"30",X"30",X"30",X"00",X"20",
		X"33",X"30",X"30",X"30",X"30",X"20",X"54",X"4F",X"20",X"20",X"35",X"30",X"30",X"30",X"30",X"00",
		X"20",X"35",X"30",X"30",X"30",X"30",X"20",X"54",X"4F",X"20",X"20",X"37",X"35",X"30",X"30",X"30",
		X"00",X"20",X"37",X"35",X"30",X"30",X"30",X"20",X"54",X"4F",X"20",X"31",X"30",X"30",X"30",X"30",
		X"30",X"00",X"20",X"20",X"20",X"20",X"20",X"4F",X"56",X"45",X"52",X"20",X"31",X"30",X"30",X"30",
		X"30",X"30",X"00",X"A9",X"E8",X"E9",X"E8",X"29",X"E9",X"69",X"E9",X"A9",X"E9",X"E9",X"E9",X"29",
		X"EA",X"69",X"EA",X"A9",X"EA",X"E9",X"EA",X"CD",X"67",X"09",X"CD",X"4C",X"09",X"CD",X"3A",X"3D",
		X"0E",X"02",X"CD",X"4E",X"3D",X"21",X"33",X"AE",X"22",X"00",X"F1",X"AF",X"32",X"03",X"F1",X"CD",
		X"C3",X"A3",X"DD",X"2A",X"00",X"F1",X"DD",X"7E",X"07",X"32",X"06",X"F8",X"0E",X"07",X"CD",X"4E",
		X"3D",X"3A",X"03",X"F1",X"FE",X"06",X"30",X"D8",X"CD",X"EC",X"A3",X"06",X"0E",X"CD",X"F9",X"3C",
		X"DB",X"00",X"E6",X"80",X"C0",X"C5",X"CD",X"AB",X"A3",X"C1",X"C0",X"10",X"F0",X"21",X"03",X"F1",
		X"34",X"18",X"DE",X"47",X"AE",X"3B",X"AE",X"00",X"00",X"06",X"34",X"28",X"24",X"28",X"34",X"28",
		X"44",X"28",X"54",X"28",X"64",X"28",X"74",X"77",X"E8",X"6D",X"AE",X"B7",X"E8",X"7A",X"AE",X"F7",
		X"E8",X"84",X"AE",X"37",X"E9",X"8E",X"AE",X"77",X"E9",X"98",X"AE",X"B7",X"E9",X"A2",X"AE",X"F7",
		X"E9",X"AC",X"AE",X"7A",X"EA",X"B6",X"AE",X"BA",X"EA",X"CF",X"AE",X"00",X"00",X"43",X"48",X"41",
		X"4E",X"4E",X"45",X"4C",X"20",X"54",X"45",X"53",X"54",X"00",X"43",X"48",X"41",X"4E",X"4E",X"45",
		X"4C",X"20",X"31",X"00",X"43",X"48",X"41",X"4E",X"4E",X"45",X"4C",X"20",X"32",X"00",X"43",X"48",
		X"41",X"4E",X"4E",X"45",X"4C",X"20",X"33",X"00",X"43",X"48",X"41",X"4E",X"4E",X"45",X"4C",X"20",
		X"34",X"00",X"43",X"48",X"41",X"4E",X"4E",X"45",X"4C",X"20",X"35",X"00",X"43",X"48",X"41",X"4E",
		X"4E",X"45",X"4C",X"20",X"36",X"00",X"50",X"52",X"45",X"53",X"53",X"20",X"57",X"45",X"41",X"50",
		X"4F",X"4E",X"53",X"20",X"56",X"41",X"4E",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"54",
		X"4F",X"20",X"45",X"58",X"49",X"54",X"20",X"54",X"45",X"53",X"54",X"00",X"21",X"24",X"AF",X"22",
		X"00",X"F1",X"3E",X"08",X"AF",X"32",X"03",X"F1",X"32",X"05",X"F1",X"CD",X"67",X"09",X"CD",X"4C",
		X"09",X"CD",X"3A",X"3D",X"0E",X"02",X"CD",X"4E",X"3D",X"CD",X"C3",X"A3",X"DD",X"2A",X"00",X"F1",
		X"DD",X"7E",X"07",X"32",X"06",X"F8",X"3A",X"05",X"F1",X"B7",X"C0",X"DB",X"00",X"2F",X"E6",X"80",
		X"C8",X"CD",X"F9",X"3C",X"CD",X"77",X"A3",X"CD",X"EC",X"A3",X"CD",X"AB",X"A3",X"28",X"E7",X"CD",
		X"11",X"A4",X"18",X"C7",X"34",X"AF",X"2C",X"AF",X"C4",X"AF",X"04",X"34",X"18",X"3E",X"18",X"4E",
		X"18",X"5E",X"18",X"6E",X"98",X"E8",X"5A",X"AF",X"1A",X"E9",X"70",X"AF",X"5A",X"E9",X"8A",X"AF",
		X"9A",X"E9",X"A2",X"AF",X"DA",X"E9",X"BD",X"AF",X"5B",X"EA",X"29",X"A5",X"9B",X"EA",X"43",X"A5",
		X"FB",X"EA",X"5F",X"A5",X"3B",X"EB",X"7A",X"A5",X"00",X"00",X"53",X"45",X"4C",X"45",X"43",X"54",
		X"20",X"41",X"20",X"54",X"45",X"53",X"54",X"20",X"4F",X"52",X"20",X"45",X"58",X"49",X"54",X"00",
		X"31",X"20",X"53",X"54",X"45",X"45",X"52",X"20",X"57",X"48",X"45",X"45",X"4C",X"20",X"43",X"41",
		X"4C",X"49",X"42",X"52",X"41",X"54",X"49",X"4F",X"4E",X"00",X"32",X"20",X"47",X"41",X"53",X"20",
		X"50",X"45",X"44",X"41",X"4C",X"20",X"43",X"41",X"4C",X"49",X"42",X"52",X"41",X"54",X"49",X"4F",
		X"4E",X"00",X"33",X"20",X"4F",X"55",X"54",X"50",X"55",X"54",X"20",X"50",X"4F",X"52",X"54",X"20",
		X"56",X"45",X"52",X"49",X"46",X"49",X"43",X"41",X"54",X"49",X"4F",X"4E",X"00",X"34",X"20",X"45",
		X"58",X"49",X"54",X"00",X"CC",X"AF",X"B4",X"B1",X"A3",X"B0",X"5A",X"A6",X"CD",X"67",X"09",X"CD",
		X"4C",X"09",X"CD",X"3A",X"3D",X"DD",X"21",X"FF",X"AF",X"CD",X"D0",X"A3",X"AF",X"32",X"37",X"F4",
		X"CD",X"F9",X"3C",X"3A",X"A2",X"F0",X"21",X"0F",X"EB",X"CD",X"81",X"B2",X"CD",X"AB",X"A3",X"28",
		X"EF",X"3A",X"A2",X"F0",X"32",X"37",X"F4",X"06",X"32",X"CD",X"F9",X"3C",X"10",X"FB",X"C9",X"75",
		X"E8",X"1D",X"B0",X"B4",X"E8",X"2C",X"B0",X"5B",X"E9",X"38",X"B0",X"BB",X"E9",X"50",X"B0",X"FB",
		X"E9",X"69",X"B0",X"5B",X"EA",X"7E",X"B0",X"D5",X"EA",X"97",X"B0",X"00",X"00",X"53",X"54",X"45",
		X"45",X"52",X"49",X"4E",X"47",X"20",X"57",X"48",X"45",X"45",X"4C",X"00",X"43",X"41",X"4C",X"49",
		X"42",X"52",X"41",X"54",X"49",X"4F",X"4E",X"00",X"31",X"20",X"43",X"45",X"4E",X"54",X"45",X"52",
		X"20",X"53",X"54",X"45",X"45",X"52",X"49",X"4E",X"47",X"20",X"57",X"48",X"45",X"45",X"4C",X"00",
		X"32",X"20",X"54",X"48",X"45",X"20",X"56",X"41",X"4C",X"55",X"45",X"20",X"4F",X"46",X"20",X"54",
		X"48",X"45",X"20",X"57",X"48",X"45",X"45",X"4C",X"00",X"20",X"20",X"53",X"48",X"4F",X"55",X"4C",
		X"44",X"20",X"42",X"45",X"20",X"20",X"38",X"43",X"20",X"20",X"48",X"45",X"58",X"00",X"33",X"20",
		X"50",X"55",X"53",X"48",X"20",X"57",X"45",X"41",X"50",X"4F",X"4E",X"20",X"56",X"41",X"4E",X"20",
		X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"57",X"48",X"45",X"45",X"4C",X"20",X"56",X"41",X"4C",
		X"55",X"45",X"00",X"CD",X"67",X"09",X"CD",X"4C",X"09",X"CD",X"3A",X"3D",X"DD",X"21",X"DF",X"B0",
		X"CD",X"D0",X"A3",X"AF",X"D3",X"04",X"21",X"2E",X"EB",X"CD",X"81",X"B2",X"06",X"20",X"CD",X"F9",
		X"3C",X"10",X"FB",X"16",X"55",X"7A",X"D3",X"04",X"21",X"2E",X"EB",X"CD",X"81",X"B2",X"0E",X"80",
		X"CD",X"AB",X"A3",X"C0",X"CD",X"F9",X"3C",X"0D",X"20",X"F6",X"7A",X"2F",X"57",X"18",X"E6",X"7A",
		X"E8",X"01",X"B1",X"1B",X"E9",X"1A",X"B1",X"5B",X"E9",X"34",X"B1",X"BB",X"E9",X"4E",X"B1",X"FB",
		X"E9",X"6A",X"B1",X"5B",X"EA",X"85",X"B1",X"9B",X"EA",X"9C",X"B1",X"F3",X"EA",X"A9",X"B1",X"00",
		X"00",X"4F",X"55",X"54",X"50",X"55",X"54",X"20",X"50",X"4F",X"52",X"54",X"20",X"56",X"45",X"52",
		X"49",X"46",X"49",X"43",X"41",X"54",X"49",X"4F",X"4E",X"00",X"54",X"48",X"45",X"20",X"56",X"41",
		X"4C",X"55",X"45",X"20",X"44",X"49",X"53",X"50",X"4C",X"41",X"59",X"45",X"44",X"20",X"42",X"45",
		X"4C",X"4F",X"57",X"00",X"48",X"41",X"53",X"20",X"42",X"45",X"45",X"4E",X"20",X"4C",X"4F",X"41",
		X"44",X"45",X"44",X"20",X"49",X"4E",X"20",X"50",X"4F",X"52",X"54",X"20",X"34",X"00",X"4F",X"55",
		X"54",X"50",X"55",X"54",X"20",X"44",X"41",X"54",X"41",X"20",X"43",X"41",X"4E",X"20",X"42",X"45",
		X"20",X"56",X"45",X"52",X"49",X"46",X"49",X"45",X"44",X"00",X"55",X"53",X"49",X"4E",X"47",X"20",
		X"54",X"48",X"45",X"20",X"55",X"4E",X"49",X"56",X"45",X"52",X"53",X"41",X"4C",X"20",X"54",X"45",
		X"53",X"54",X"45",X"52",X"00",X"50",X"55",X"53",X"48",X"20",X"57",X"45",X"41",X"50",X"4F",X"4E",
		X"20",X"56",X"41",X"4E",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"54",X"4F",X"20",X"45",
		X"58",X"49",X"54",X"20",X"54",X"45",X"53",X"54",X"00",X"54",X"45",X"53",X"54",X"20",X"56",X"41",
		X"4C",X"55",X"45",X"00",X"CD",X"67",X"09",X"CD",X"4C",X"09",X"CD",X"3A",X"3D",X"DD",X"21",X"EB",
		X"B1",X"CD",X"D0",X"A3",X"AF",X"32",X"38",X"F4",X"CD",X"F9",X"3C",X"3A",X"7E",X"F0",X"C6",X"02",
		X"21",X"0F",X"EB",X"CD",X"81",X"B2",X"CD",X"AB",X"A3",X"28",X"ED",X"3A",X"7E",X"F0",X"C6",X"02",
		X"32",X"38",X"F4",X"06",X"32",X"CD",X"F9",X"3C",X"10",X"FB",X"C9",X"75",X"E8",X"09",X"B2",X"B5",
		X"E8",X"13",X"B2",X"5B",X"E9",X"1F",X"B2",X"BB",X"E9",X"33",X"B2",X"FB",X"E9",X"49",X"B2",X"5B",
		X"EA",X"58",X"B2",X"D6",X"EA",X"71",X"B2",X"00",X"00",X"47",X"41",X"53",X"20",X"50",X"45",X"44",
		X"41",X"4C",X"00",X"43",X"41",X"4C",X"49",X"42",X"52",X"41",X"54",X"49",X"4F",X"4E",X"00",X"31",
		X"20",X"52",X"45",X"4C",X"45",X"41",X"53",X"45",X"20",X"47",X"41",X"53",X"20",X"50",X"45",X"44",
		X"41",X"4C",X"00",X"32",X"20",X"54",X"48",X"45",X"20",X"47",X"41",X"53",X"20",X"50",X"45",X"44",
		X"41",X"4C",X"20",X"56",X"41",X"4C",X"55",X"45",X"00",X"20",X"20",X"53",X"48",X"4F",X"55",X"4C",
		X"44",X"20",X"42",X"45",X"20",X"30",X"42",X"00",X"33",X"20",X"50",X"55",X"53",X"48",X"20",X"57",
		X"45",X"41",X"50",X"4F",X"4E",X"20",X"56",X"41",X"4E",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",
		X"00",X"47",X"41",X"53",X"20",X"50",X"45",X"44",X"41",X"4C",X"20",X"56",X"41",X"4C",X"55",X"45",
		X"00",X"C5",X"47",X"0E",X"02",X"E6",X"0F",X"C6",X"30",X"FE",X"3A",X"38",X"02",X"C6",X"07",X"BE",
		X"28",X"01",X"77",X"78",X"0D",X"28",X"0A",X"23",X"78",X"06",X"00",X"0F",X"0F",X"0F",X"0F",X"18",
		X"E4",X"C1",X"C9",X"CD",X"67",X"09",X"CD",X"4C",X"09",X"CD",X"3A",X"3D",X"0E",X"02",X"CD",X"4E",
		X"3D",X"DD",X"21",X"CA",X"B2",X"CD",X"D0",X"A3",X"AF",X"32",X"09",X"F1",X"DB",X"00",X"2F",X"E6",
		X"80",X"C8",X"CD",X"F9",X"3C",X"CD",X"45",X"B3",X"18",X"F2",X"76",X"E8",X"DC",X"B2",X"1A",X"EB",
		X"EA",X"B2",X"3A",X"EB",X"04",X"B3",X"7A",X"EB",X"19",X"B3",X"00",X"00",X"50",X"4C",X"41",X"59",
		X"45",X"52",X"20",X"49",X"4E",X"50",X"55",X"54",X"53",X"00",X"41",X"43",X"54",X"49",X"56",X"41",
		X"54",X"45",X"20",X"41",X"4C",X"4C",X"20",X"50",X"4C",X"41",X"59",X"45",X"52",X"20",X"49",X"4E",
		X"50",X"55",X"54",X"00",X"53",X"57",X"49",X"54",X"43",X"48",X"45",X"53",X"20",X"41",X"4E",X"44",
		X"20",X"44",X"45",X"56",X"49",X"43",X"45",X"53",X"00",X"48",X"49",X"54",X"20",X"54",X"49",X"4C",
		X"54",X"20",X"54",X"4F",X"20",X"45",X"58",X"49",X"54",X"00",X"43",X"45",X"4E",X"54",X"45",X"52",
		X"45",X"44",X"00",X"52",X"49",X"47",X"48",X"54",X"20",X"20",X"20",X"00",X"4C",X"45",X"46",X"54",
		X"20",X"20",X"20",X"20",X"00",X"DD",X"21",X"58",X"B4",X"FD",X"21",X"0A",X"F1",X"DD",X"7E",X"00",
		X"FE",X"FF",X"CA",X"54",X"B4",X"B7",X"CA",X"5F",X"B3",X"F2",X"D8",X"B3",X"C3",X"4A",X"B4",X"06",
		X"00",X"DD",X"4E",X"01",X"ED",X"78",X"2F",X"DD",X"A6",X"02",X"47",X"FD",X"BE",X"00",X"20",X"07",
		X"3A",X"09",X"F1",X"B7",X"C2",X"4A",X"B4",X"FD",X"70",X"00",X"78",X"DD",X"6E",X"04",X"DD",X"66",
		X"05",X"4E",X"23",X"46",X"23",X"B7",X"28",X"27",X"3A",X"12",X"F0",X"DD",X"B6",X"08",X"32",X"12",
		X"F0",X"EB",X"C5",X"E1",X"CD",X"18",X"3F",X"3A",X"09",X"F1",X"B7",X"CA",X"4A",X"B4",X"0E",X"02",
		X"CD",X"4E",X"3D",X"CD",X"F9",X"3C",X"DD",X"4E",X"03",X"CD",X"4E",X"3D",X"C3",X"4A",X"B4",X"3A",
		X"09",X"F1",X"B7",X"28",X"0B",X"3A",X"12",X"F0",X"DD",X"AE",X"08",X"32",X"12",X"F0",X"18",X"0B",
		X"32",X"12",X"F0",X"3A",X"5C",X"F0",X"F6",X"04",X"32",X"5C",X"F0",X"DD",X"5E",X"06",X"DD",X"56",
		X"07",X"C5",X"E1",X"CD",X"18",X"3F",X"18",X"72",X"3A",X"09",X"F1",X"B7",X"20",X"10",X"DD",X"6E",
		X"04",X"DD",X"66",X"05",X"4E",X"23",X"46",X"23",X"EB",X"C5",X"E1",X"CD",X"18",X"3F",X"DD",X"7E",
		X"00",X"FE",X"01",X"20",X"3B",X"3A",X"A1",X"F0",X"FD",X"BE",X"00",X"20",X"09",X"3A",X"C8",X"E8",
		X"B7",X"20",X"47",X"3A",X"A1",X"F0",X"FD",X"77",X"00",X"21",X"C9",X"E8",X"B7",X"28",X"19",X"CB",
		X"7F",X"11",X"3C",X"B3",X"28",X"05",X"11",X"33",X"B3",X"ED",X"44",X"F5",X"CD",X"18",X"3F",X"F1",
		X"F6",X"30",X"21",X"C3",X"E8",X"77",X"18",X"22",X"11",X"2A",X"B3",X"CD",X"18",X"3F",X"18",X"1A",
		X"3A",X"7E",X"F0",X"FD",X"BE",X"00",X"20",X"09",X"3A",X"E8",X"E8",X"B7",X"20",X"0C",X"3A",X"7E",
		X"F0",X"FD",X"77",X"00",X"21",X"E8",X"E8",X"CD",X"81",X"B2",X"11",X"09",X"00",X"DD",X"19",X"FD",
		X"23",X"C3",X"4D",X"B3",X"32",X"09",X"F1",X"C9",X"01",X"02",X"FF",X"01",X"CE",X"B4",X"CE",X"B4",
		X"00",X"02",X"02",X"FF",X"01",X"E1",X"B4",X"E1",X"B4",X"00",X"00",X"00",X"10",X"01",X"EF",X"B4",
		X"01",X"B5",X"00",X"00",X"01",X"10",X"37",X"2F",X"B5",X"E8",X"B5",X"01",X"00",X"01",X"01",X"24",
		X"3E",X"B5",X"E8",X"B5",X"08",X"00",X"01",X"08",X"25",X"4C",X"B5",X"E8",X"B5",X"02",X"00",X"00",
		X"01",X"0C",X"5B",X"B5",X"E8",X"B5",X"00",X"00",X"00",X"02",X"0C",X"6A",X"B5",X"E8",X"B5",X"00",
		X"00",X"00",X"40",X"0B",X"79",X"B5",X"E8",X"B5",X"00",X"00",X"01",X"02",X"30",X"20",X"B5",X"E8",
		X"B5",X"80",X"00",X"01",X"04",X"4F",X"11",X"B5",X"E8",X"B5",X"04",X"00",X"03",X"02",X"01",X"8A",
		X"B5",X"A1",X"B5",X"00",X"00",X"03",X"01",X"01",X"B6",X"B5",X"D0",X"B5",X"00",X"FF",X"D9",X"E8",
		X"53",X"54",X"45",X"45",X"52",X"49",X"4E",X"47",X"20",X"57",X"48",X"45",X"45",X"4C",X"20",X"20",
		X"00",X"F9",X"E8",X"47",X"41",X"53",X"20",X"50",X"45",X"44",X"41",X"4C",X"20",X"20",X"00",X"19",
		X"E9",X"47",X"45",X"41",X"52",X"20",X"53",X"48",X"49",X"46",X"54",X"20",X"48",X"49",X"47",X"48",
		X"00",X"47",X"45",X"41",X"52",X"20",X"53",X"48",X"49",X"46",X"54",X"20",X"4C",X"4F",X"57",X"20",
		X"00",X"39",X"E9",X"57",X"45",X"41",X"50",X"4F",X"4E",X"20",X"54",X"52",X"55",X"43",X"4B",X"00",
		X"59",X"E9",X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"53",X"20",X"20",X"20",X"20",X"00",X"79",
		X"E9",X"4D",X"41",X"43",X"48",X"49",X"4E",X"45",X"20",X"47",X"55",X"4E",X"20",X"00",X"99",X"E9",
		X"4F",X"49",X"4C",X"20",X"53",X"4C",X"49",X"43",X"4B",X"20",X"20",X"00",X"B9",X"E9",X"53",X"4D",
		X"4F",X"4B",X"45",X"20",X"53",X"43",X"52",X"45",X"45",X"4E",X"00",X"F9",X"E9",X"43",X"4F",X"49",
		X"4E",X"20",X"43",X"48",X"55",X"54",X"45",X"20",X"31",X"00",X"19",X"EA",X"43",X"4F",X"49",X"4E",
		X"20",X"43",X"48",X"55",X"54",X"45",X"20",X"32",X"00",X"39",X"EA",X"53",X"45",X"52",X"56",X"49",
		X"43",X"45",X"20",X"42",X"55",X"54",X"54",X"4F",X"4E",X"00",X"79",X"EA",X"4D",X"55",X"53",X"49",
		X"43",X"20",X"49",X"4E",X"20",X"41",X"54",X"54",X"52",X"41",X"43",X"54",X"20",X"53",X"45",X"51",
		X"00",X"53",X"49",X"4C",X"45",X"4E",X"54",X"20",X"41",X"54",X"54",X"52",X"41",X"43",X"54",X"20",
		X"53",X"45",X"51",X"20",X"20",X"00",X"B9",X"EA",X"31",X"20",X"4D",X"49",X"4E",X"55",X"54",X"45",
		X"20",X"47",X"41",X"4D",X"45",X"20",X"54",X"49",X"4D",X"45",X"52",X"20",X"20",X"20",X"20",X"00",
		X"31",X"20",X"4D",X"49",X"4E",X"20",X"33",X"30",X"20",X"53",X"45",X"43",X"20",X"47",X"41",X"4D",
		X"45",X"20",X"54",X"49",X"4D",X"45",X"52",X"00",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",
		X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"20",X"00",X"CD",X"67",X"09",X"CD",X"4C",X"09",
		X"CD",X"3A",X"3D",X"DD",X"21",X"51",X"B7",X"CD",X"D0",X"A3",X"DD",X"21",X"7E",X"B8",X"DD",X"7E",
		X"00",X"FE",X"BF",X"28",X"0A",X"CD",X"1A",X"B7",X"11",X"06",X"00",X"DD",X"19",X"18",X"EF",X"FD",
		X"21",X"04",X"F8",X"FD",X"36",X"00",X"28",X"FD",X"36",X"02",X"34",X"DD",X"21",X"7E",X"B8",X"DD",
		X"7E",X"00",X"FD",X"77",X"03",X"DB",X"00",X"E6",X"80",X"C0",X"DB",X"01",X"2F",X"E6",X"08",X"20",
		X"1B",X"DB",X"01",X"2F",X"E6",X"01",X"28",X"35",X"DD",X"7E",X"00",X"FE",X"BF",X"28",X"07",X"01",
		X"06",X"00",X"DD",X"09",X"18",X"1D",X"DD",X"21",X"7E",X"B8",X"18",X"17",X"DD",X"7E",X"00",X"FE",
		X"27",X"28",X"07",X"01",X"FA",X"FF",X"DD",X"09",X"18",X"09",X"DD",X"21",X"A8",X"B8",X"18",X"03",
		X"DD",X"7E",X"00",X"DD",X"7E",X"00",X"FD",X"77",X"03",X"AF",X"32",X"0A",X"F1",X"DB",X"01",X"E6",
		X"02",X"20",X"27",X"DD",X"7E",X"00",X"FE",X"BF",X"C8",X"DD",X"6E",X"02",X"DD",X"66",X"03",X"7E",
		X"FE",X"09",X"30",X"03",X"34",X"18",X"62",X"DD",X"7E",X"01",X"FE",X"01",X"28",X"0C",X"2B",X"7E",
		X"FE",X"09",X"28",X"06",X"34",X"23",X"36",X"00",X"18",X"4F",X"DB",X"01",X"E6",X"10",X"28",X"06",
		X"AF",X"32",X"0A",X"F1",X"18",X"51",X"DD",X"7E",X"00",X"FE",X"BF",X"C8",X"DD",X"6E",X"02",X"DD",
		X"66",X"03",X"7E",X"FE",X"02",X"38",X"03",X"35",X"18",X"2F",X"DD",X"7E",X"01",X"FE",X"01",X"28",
		X"36",X"7E",X"B7",X"20",X"1D",X"36",X"09",X"2B",X"35",X"7E",X"FE",X"01",X"20",X"1B",X"D5",X"11",
		X"33",X"F4",X"7D",X"BB",X"20",X"09",X"7C",X"BA",X"20",X"05",X"36",X"02",X"23",X"36",X"00",X"D1",
		X"18",X"07",X"2B",X"7E",X"B7",X"28",X"10",X"23",X"35",X"CD",X"1A",X"B7",X"3A",X"0A",X"F1",X"FE",
		X"04",X"30",X"04",X"3C",X"32",X"0A",X"F1",X"3A",X"0A",X"F1",X"06",X"06",X"FE",X"03",X"38",X"02",
		X"06",X"01",X"CD",X"F9",X"3C",X"10",X"FB",X"C3",X"35",X"B6",X"DD",X"46",X"01",X"21",X"19",X"F1",
		X"DD",X"5E",X"02",X"DD",X"56",X"03",X"78",X"3D",X"28",X"01",X"1B",X"1A",X"B7",X"20",X"08",X"78",
		X"3D",X"28",X"04",X"3E",X"20",X"18",X"02",X"C6",X"30",X"77",X"23",X"13",X"10",X"ED",X"36",X"00",
		X"11",X"19",X"F1",X"DD",X"4E",X"04",X"DD",X"46",X"05",X"C5",X"E1",X"CD",X"18",X"3F",X"C3",X"F9",
		X"3C",X"55",X"E8",X"A3",X"B7",X"9A",X"E8",X"C9",X"B7",X"8F",X"E8",X"B1",X"B7",X"B3",X"E8",X"74",
		X"B8",X"D3",X"E8",X"C1",X"B7",X"1A",X"E9",X"C9",X"B7",X"0F",X"E9",X"B3",X"B7",X"33",X"E9",X"74",
		X"B8",X"53",X"E9",X"C1",X"B7",X"9A",X"E9",X"28",X"B8",X"FA",X"E9",X"D4",X"B7",X"15",X"EA",X"EE",
		X"B7",X"5A",X"EA",X"FA",X"B7",X"75",X"EA",X"EE",X"B7",X"96",X"EA",X"13",X"B8",X"16",X"EB",X"39",
		X"B8",X"5B",X"EB",X"29",X"A5",X"7B",X"EB",X"43",X"A5",X"BB",X"EB",X"3E",X"B8",X"DB",X"EB",X"5A",
		X"B8",X"00",X"00",X"53",X"45",X"54",X"55",X"50",X"20",X"4F",X"50",X"54",X"49",X"4F",X"4E",X"53",
		X"00",X"31",X"00",X"32",X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"20",X"46",X"4F",X"52",
		X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"00",X"43",X"4F",X"49",X"4E",X"20",X"43",X"48",
		X"55",X"54",X"45",X"00",X"31",X"53",X"54",X"20",X"45",X"58",X"54",X"52",X"41",X"20",X"42",X"41",
		X"53",X"45",X"20",X"41",X"57",X"41",X"52",X"44",X"45",X"44",X"20",X"41",X"54",X"00",X"30",X"30",
		X"30",X"30",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",X"00",X"45",X"58",X"54",X"52",X"41",X"20",
		X"42",X"41",X"53",X"45",X"20",X"41",X"57",X"41",X"52",X"44",X"45",X"44",X"20",X"45",X"56",X"45",
		X"52",X"59",X"00",X"55",X"50",X"20",X"54",X"4F",X"20",X"41",X"20",X"4D",X"41",X"58",X"49",X"4D",
		X"55",X"4D",X"20",X"4F",X"46",X"20",X"33",X"00",X"44",X"49",X"46",X"46",X"49",X"43",X"55",X"4C",
		X"54",X"59",X"20",X"4C",X"45",X"56",X"45",X"4C",X"00",X"45",X"58",X"49",X"54",X"00",X"55",X"53",
		X"45",X"20",X"4D",X"49",X"53",X"53",X"49",X"4C",X"45",X"20",X"41",X"4E",X"44",X"20",X"4D",X"41",
		X"43",X"48",X"49",X"4E",X"45",X"20",X"47",X"55",X"4E",X"00",X"54",X"52",X"49",X"47",X"47",X"45",
		X"52",X"53",X"20",X"54",X"4F",X"20",X"43",X"48",X"41",X"4E",X"47",X"45",X"20",X"56",X"41",X"4C",
		X"55",X"45",X"53",X"00",X"43",X"4F",X"49",X"4E",X"53",X"20",X"46",X"4F",X"52",X"00",X"27",X"01",
		X"2B",X"F4",X"B6",X"E8",X"2F",X"01",X"2C",X"F4",X"D6",X"E8",X"47",X"01",X"2D",X"F4",X"36",X"E9",
		X"4F",X"01",X"2E",X"F4",X"56",X"E9",X"67",X"01",X"32",X"F4",X"B6",X"E9",X"7F",X"02",X"34",X"F4",
		X"16",X"EA",X"97",X"02",X"36",X"F4",X"76",X"EA",X"BF",X"54",X"4F",X"20",X"53",X"54",X"41",X"52",
		X"54",X"00",X"50",X"52",X"45",X"53",X"53",X"20",X"54",X"48",X"45",X"20",X"46",X"4C",X"41",X"53",
		X"48",X"49",X"4E",X"47",X"00",X"53",X"54",X"45",X"45",X"52",X"49",X"4E",X"47",X"20",X"57",X"48",
		X"45",X"45",X"4C",X"20",X"48",X"55",X"42",X"00",X"4F",X"52",X"20",X"50",X"52",X"45",X"53",X"53",
		X"00",X"41",X"43",X"43",X"45",X"4C",X"45",X"52",X"41",X"54",X"4F",X"52",X"20",X"20",X"50",X"45",
		X"44",X"41",X"4C",X"00",X"20",X"46",X"4F",X"52",X"20",X"49",X"4E",X"53",X"54",X"52",X"55",X"43",
		X"54",X"49",X"4F",X"4E",X"53",X"20",X"00",X"49",X"4E",X"53",X"45",X"52",X"54",X"20",X"20",X"43",
		X"4F",X"49",X"4E",X"00",X"43",X"52",X"45",X"44",X"49",X"54",X"53",X"00",X"47",X"41",X"4D",X"45",
		X"20",X"20",X"4F",X"56",X"45",X"52",X"00",X"49",X"43",X"59",X"00",X"52",X"4F",X"41",X"44",X"53",
		X"00",X"41",X"48",X"45",X"41",X"44",X"00",X"4E",X"4F",X"20",X"50",X"4F",X"49",X"4E",X"54",X"53",
		X"00",X"48",X"49",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"00",X"00",X"00",X"00",
		X"02",X"05",X"00",X"00",X"00",X"00",X"01",X"05",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"00",X"00",X"1A",X"00",X"00",X"00",X"00",X"10",X"1C",X"00",X"0A",
		X"02",X"FA",X"02",X"1C",X"10",X"0A",X"02",X"FA",X"02",X"1A",X"10",X"00",X"04",X"00",X"F4",X"1A",
		X"30",X"00",X"04",X"00",X"F4",X"1C",X"30",X"F6",X"02",X"06",X"02",X"1C",X"20",X"F6",X"02",X"06",
		X"02",X"1A",X"20",X"00",X"00",X"00",X"10",X"21",X"00",X"00",X"00",X"00",X"10",X"84",X"00",X"00",
		X"00",X"00",X"10",X"84",X"00",X"00",X"00",X"00",X"10",X"84",X"00",X"00",X"00",X"00",X"10",X"84",
		X"00",X"00",X"00",X"00",X"10",X"84",X"00",X"00",X"00",X"00",X"10",X"84",X"00",X"00",X"00",X"00",
		X"10",X"84",X"00",X"00",X"00",X"00",X"10",X"84",X"00",X"00",X"00",X"00",X"10",X"84",X"00",X"00",
		X"00",X"00",X"10",X"D4",X"00",X"00",X"00",X"00",X"10",X"03",X"06",X"23",X"14",X"06",X"2C",X"02",
		X"06",X"24",X"03",X"07",X"23",X"14",X"07",X"2C",X"11",X"08",X"27",X"03",X"08",X"23",X"02",X"09",
		X"24",X"11",X"09",X"27",X"10",X"00",X"25",X"00",X"00",X"00",X"71",X"FF",X"27",X"11",X"0C",X"7C",
		X"14",X"06",X"2C",X"02",X"06",X"24",X"71",X"0C",X"27",X"03",X"05",X"23",X"14",X"07",X"2C",X"71",
		X"0D",X"27",X"02",X"09",X"24",X"10",X"00",X"25",X"16",X"6A",X"00",X"71",X"FF",X"27",X"11",X"0C",
		X"7C",X"14",X"06",X"2C",X"02",X"06",X"24",X"71",X"0A",X"27",X"03",X"07",X"23",X"11",X"0B",X"7C",
		X"03",X"08",X"23",X"71",X"0C",X"27",X"10",X"00",X"25",X"17",X"6B",X"00",X"71",X"FF",X"27",X"11",
		X"0A",X"7C",X"03",X"06",X"23",X"14",X"04",X"2C",X"71",X"0C",X"27",X"03",X"05",X"23",X"71",X"09",
		X"27",X"14",X"07",X"2C",X"11",X"0C",X"7C",X"10",X"00",X"25",X"17",X"6B",X"00",X"71",X"FF",X"27",
		X"11",X"0C",X"7C",X"71",X"0A",X"27",X"14",X"06",X"2C",X"11",X"0C",X"7C",X"02",X"09",X"24",X"71",
		X"0D",X"27",X"03",X"08",X"23",X"11",X"0C",X"7C",X"10",X"00",X"25",X"18",X"69",X"00",X"71",X"FF",
		X"27",X"11",X"0B",X"7C",X"71",X"0C",X"27",X"14",X"06",X"2C",X"11",X"0B",X"7C",X"14",X"07",X"2C",
		X"02",X"08",X"24",X"71",X"0D",X"27",X"03",X"08",X"23",X"10",X"00",X"25",X"16",X"6A",X"00",X"71",
		X"FF",X"27",X"11",X"0C",X"7C",X"71",X"0D",X"27",X"14",X"06",X"2C",X"11",X"0C",X"7C",X"02",X"09",
		X"24",X"71",X"0D",X"27",X"03",X"08",X"23",X"11",X"0C",X"7C",X"10",X"00",X"25",X"16",X"6A",X"00",
		X"91",X"09",X"70",X"91",X"08",X"70",X"91",X"08",X"70",X"91",X"09",X"70",X"91",X"07",X"70",X"91",
		X"0A",X"70",X"91",X"06",X"70",X"91",X"07",X"70",X"91",X"0B",X"70",X"90",X"00",X"AB",X"00",X"00",
		X"00",X"20",X"14",X"10",X"10",X"14",X"20",X"28",X"28",X"28",X"06",X"04",X"01",X"02",X"04",X"07",
		X"07",X"07",X"07",X"05",X"BB",X"0D",X"BB",X"15",X"BB",X"1D",X"BB",X"25",X"BB",X"2D",X"BB",X"35",
		X"BB",X"3D",X"BB",X"45",X"BB",X"01",X"02",X"03",X"03",X"04",X"04",X"05",X"05",X"02",X"03",X"03",
		X"04",X"04",X"05",X"05",X"06",X"02",X"03",X"04",X"04",X"05",X"05",X"06",X"06",X"03",X"04",X"04",
		X"05",X"05",X"06",X"06",X"06",X"03",X"04",X"05",X"05",X"05",X"06",X"06",X"06",X"03",X"04",X"05",
		X"05",X"06",X"06",X"06",X"06",X"03",X"04",X"05",X"06",X"06",X"06",X"06",X"06",X"04",X"05",X"05",
		X"06",X"06",X"06",X"06",X"06",X"04",X"05",X"06",X"06",X"06",X"06",X"06",X"06",X"00",X"00",X"00",
		X"00",X"04",X"06",X"04",X"08",X"06",X"06",X"04",X"08",X"00",X"10",X"00",X"10",X"02",X"0C",X"02",
		X"0C",X"06",X"04",X"06",X"04",X"02",X"0C",X"00",X"0C",X"04",X"08",X"06",X"04",X"00",X"10",X"00",
		X"10",X"0A",X"09",X"F8",X"FA",X"00",X"F8",X"F8",X"3F",X"F8",X"32",X"0C",X"07",X"F6",X"FC",X"10",
		X"F6",X"FC",X"17",X"F1",X"6D",X"07",X"05",X"F9",X"01",X"10",X"E9",X"02",X"14",X"E8",X"6D",X"08",
		X"03",X"FA",X"08",X"10",X"EA",X"0D",X"3E",X"E8",X"31",X"08",X"05",X"F9",X"0E",X"30",X"E9",X"11",
		X"14",X"EA",X"33",X"04",X"07",X"F6",X"14",X"30",X"F6",X"16",X"17",X"F5",X"33",X"06",X"09",X"F8",
		X"16",X"30",X"F8",X"17",X"3F",X"F8",X"32",X"04",X"07",X"FA",X"14",X"20",X"FA",X"14",X"17",X"FF",
		X"6D",X"09",X"05",X"F7",X"0F",X"20",X"07",X"0E",X"14",X"09",X"6D",X"08",X"03",X"F6",X"08",X"00",
		X"06",X"09",X"3E",X"08",X"31",X"07",X"05",X"F7",X"01",X"00",X"07",X"FE",X"14",X"06",X"33",X"0B",
		X"07",X"FA",X"FB",X"00",X"FA",X"F9",X"17",X"FB",X"33",X"08",X"51",X"F6",X"08",X"00",X"06",X"09",
		X"3E",X"07",X"31",X"FF",X"BB",X"0B",X"BC",X"17",X"BC",X"23",X"BC",X"2F",X"BC",X"3B",X"BC",X"AE",
		X"00",X"B0",X"00",X"AF",X"00",X"B1",X"00",X"B4",X"00",X"B5",X"00",X"B0",X"20",X"AE",X"20",X"B1",
		X"20",X"AF",X"20",X"B5",X"20",X"B4",X"20",X"B2",X"00",X"B0",X"00",X"B3",X"00",X"B1",X"00",X"B6",
		X"00",X"B5",X"00",X"B0",X"20",X"B2",X"20",X"B1",X"20",X"B3",X"20",X"B5",X"20",X"B6",X"20",X"AE",
		X"00",X"AE",X"20",X"AF",X"00",X"AF",X"20",X"B4",X"00",X"B4",X"20",X"B2",X"00",X"B2",X"20",X"B3",
		X"00",X"B3",X"20",X"B6",X"00",X"B6",X"20",X"23",X"C9",X"D9",X"B9",X"B1",X"BF",X"04",X"00",X"BB",
		X"BF",X"03",X"00",X"CF",X"BF",X"DD",X"BF",X"EF",X"BF",X"04",X"00",X"F9",X"BF",X"06",X"00",X"03",
		X"C0",X"0D",X"C0",X"3D",X"C0",X"F9",X"BF",X"49",X"C0",X"53",X"C0",X"06",X"00",X"53",X"C0",X"83",
		X"C0",X"EF",X"BF",X"03",X"00",X"B5",X"C0",X"DB",X"C0",X"E5",X"C0",X"07",X"00",X"2F",X"C1",X"00",
		X"00",X"85",X"BC",X"DB",X"BC",X"43",X"C9",X"FA",X"B9",X"3D",X"C1",X"49",X"C1",X"C5",X"BF",X"10",
		X"00",X"CF",X"BF",X"DD",X"BF",X"F9",X"BF",X"05",X"00",X"49",X"C0",X"53",X"C0",X"03",X"00",X"5D",
		X"C0",X"6B",X"C0",X"6B",X"C0",X"75",X"C0",X"53",X"C0",X"06",X"00",X"83",X"C0",X"03",X"C0",X"3D",
		X"C0",X"EF",X"BF",X"F9",X"BF",X"EF",X"BF",X"F9",X"BF",X"EF",X"BF",X"F9",X"BF",X"8F",X"C0",X"9D",
		X"C0",X"02",X"00",X"A7",X"C0",X"EF",X"BF",X"F9",X"BF",X"F9",X"BF",X"B5",X"C0",X"DB",X"C0",X"E5",
		X"C0",X"07",X"00",X"2F",X"C1",X"00",X"00",X"23",X"BD",X"7D",X"BD",X"63",X"C9",X"1B",X"BA",X"57",
		X"C1",X"65",X"C1",X"B1",X"BF",X"03",X"00",X"BB",X"BF",X"03",X"00",X"C5",X"BF",X"03",X"00",X"BB",
		X"BF",X"07",X"00",X"B1",X"BF",X"03",X"00",X"CF",X"BF",X"DD",X"BF",X"EF",X"BF",X"F9",X"BF",X"EF",
		X"BF",X"F9",X"BF",X"B5",X"C0",X"C5",X"BF",X"BB",X"BF",X"DB",X"C0",X"E5",X"C0",X"12",X"00",X"EF",
		X"C0",X"F9",X"C0",X"07",X"C1",X"05",X"00",X"11",X"C1",X"E5",X"C0",X"2F",X"C1",X"00",X"00",X"D9",
		X"BD",X"7D",X"BD",X"63",X"C9",X"3C",X"BA",X"3D",X"C1",X"49",X"C1",X"C5",X"BF",X"07",X"00",X"B1",
		X"BF",X"0D",X"00",X"C5",X"BF",X"03",X"00",X"CF",X"BF",X"DD",X"BF",X"EF",X"BF",X"03",X"00",X"F9",
		X"BF",X"03",X"C0",X"0D",X"C0",X"17",X"C0",X"25",X"C0",X"03",X"00",X"2F",X"C0",X"0D",X"C0",X"3D",
		X"C0",X"49",X"C0",X"53",X"C0",X"02",X"00",X"83",X"C0",X"EF",X"BF",X"03",X"00",X"EF",X"BF",X"B5",
		X"C0",X"BB",X"BF",X"DB",X"C0",X"E5",X"C0",X"04",X"00",X"EF",X"C0",X"F9",X"C0",X"07",X"C1",X"07",
		X"C1",X"11",X"C1",X"E5",X"C0",X"2F",X"C1",X"00",X"00",X"7F",X"BE",X"7D",X"BD",X"A3",X"C9",X"5D",
		X"BA",X"57",X"C1",X"65",X"C1",X"C5",X"BF",X"07",X"00",X"CF",X"BF",X"DD",X"BF",X"EF",X"BF",X"05",
		X"00",X"49",X"C0",X"53",X"C0",X"07",X"00",X"83",X"C0",X"49",X"C0",X"83",X"C0",X"03",X"C0",X"3D",
		X"C0",X"F9",X"BF",X"03",X"00",X"8F",X"C0",X"9D",X"C0",X"05",X"00",X"A7",X"C0",X"EF",X"BF",X"03",
		X"00",X"03",X"C0",X"3D",X"C0",X"49",X"C0",X"83",X"C0",X"03",X"C0",X"3D",X"C0",X"03",X"C0",X"3D",
		X"C0",X"EF",X"BF",X"B5",X"C0",X"C5",X"BF",X"BB",X"BF",X"C5",X"BF",X"DB",X"C0",X"E5",X"C0",X"06",
		X"00",X"2F",X"C1",X"00",X"00",X"7F",X"BE",X"01",X"BE",X"C3",X"C9",X"7E",X"BA",X"3D",X"C1",X"49",
		X"C1",X"B1",X"BF",X"1F",X"00",X"DB",X"C0",X"E5",X"C0",X"12",X"00",X"EF",X"C0",X"F9",X"C0",X"07",
		X"C1",X"07",X"00",X"11",X"C1",X"E5",X"C0",X"03",X"00",X"2F",X"C1",X"00",X"00",X"85",X"BC",X"01",
		X"BE",X"23",X"C9",X"9F",X"BA",X"57",X"C1",X"65",X"C1",X"B1",X"BF",X"BB",X"BF",X"03",X"00",X"C5",
		X"BF",X"03",X"00",X"CF",X"BF",X"DD",X"BF",X"EF",X"BF",X"03",X"C0",X"0D",X"C0",X"0D",X"C0",X"17",
		X"C0",X"25",X"C0",X"02",X"00",X"2F",X"C0",X"3D",X"C0",X"F9",X"BF",X"8F",X"C0",X"9D",X"C0",X"A7",
		X"C0",X"49",X"C0",X"83",X"C0",X"03",X"C0",X"3D",X"C0",X"03",X"C0",X"3D",X"C0",X"03",X"C0",X"3D",
		X"C0",X"49",X"C0",X"83",X"C0",X"49",X"C0",X"53",X"C0",X"73",X"C1",X"7F",X"C1",X"89",X"C1",X"AB",
		X"C1",X"6B",X"C0",X"00",X"01",X"6B",X"C0",X"C1",X"C1",X"CF",X"C1",X"D9",X"C1",X"53",X"C0",X"83",
		X"C0",X"EF",X"BF",X"B5",X"C0",X"BB",X"BF",X"DB",X"C0",X"E5",X"C0",X"EF",X"C0",X"F9",X"C0",X"07",
		X"C1",X"07",X"00",X"11",X"C1",X"E5",X"C0",X"2F",X"C1",X"00",X"00",X"85",X"BC",X"DB",X"BC",X"23",
		X"C9",X"5D",X"BA",X"3D",X"C1",X"49",X"C1",X"B1",X"BF",X"06",X"00",X"BB",X"BF",X"04",X"00",X"CF",
		X"BF",X"DD",X"BF",X"EF",X"BF",X"02",X"00",X"03",X"C0",X"0D",X"C0",X"03",X"00",X"3D",X"C0",X"F9",
		X"BF",X"03",X"00",X"49",X"C0",X"83",X"C0",X"03",X"C0",X"3D",X"C0",X"03",X"C0",X"3D",X"C0",X"03",
		X"C0",X"3D",X"C0",X"49",X"C0",X"83",X"C0",X"49",X"C0",X"53",X"C0",X"02",X"00",X"73",X"C1",X"7F",
		X"C1",X"89",X"C1",X"AB",X"C1",X"6B",X"C0",X"00",X"01",X"6B",X"C0",X"C1",X"C1",X"CF",X"C1",X"D9",
		X"C1",X"53",X"C0",X"83",X"C0",X"EF",X"BF",X"03",X"00",X"B5",X"C0",X"DB",X"C0",X"E5",X"C0",X"07",
		X"00",X"2F",X"C1",X"00",X"00",X"D9",X"BD",X"DB",X"BC",X"23",X"C9",X"C0",X"BA",X"97",X"C3",X"E3",
		X"C1",X"05",X"00",X"ED",X"C1",X"FF",X"C1",X"0D",X"C2",X"07",X"00",X"17",X"C2",X"29",X"C2",X"FF",
		X"C1",X"53",X"C2",X"1B",X"C3",X"F7",X"C2",X"02",X"00",X"01",X"C3",X"11",X"C3",X"29",X"C3",X"29",
		X"C2",X"1B",X"C3",X"F7",X"C2",X"01",X"C3",X"29",X"C3",X"29",X"C2",X"1B",X"C3",X"6F",X"C2",X"89",
		X"C3",X"7D",X"C2",X"97",X"C2",X"AF",X"C2",X"BD",X"C2",X"CF",X"C2",X"D9",X"C2",X"F7",X"C2",X"03",
		X"00",X"01",X"C3",X"29",X"C3",X"29",X"C2",X"3D",X"C2",X"0D",X"C2",X"05",X"00",X"00",X"00",X"67",
		X"BF",X"23",X"C9",X"5D",X"BA",X"53",X"C0",X"45",X"C3",X"4F",X"C3",X"73",X"C3",X"7D",X"C3",X"53",
		X"C0",X"83",X"C0",X"EF",X"BF",X"03",X"00",X"B5",X"C0",X"DB",X"C0",X"E5",X"C0",X"07",X"00",X"2F",
		X"C1",X"00",X"00",X"D9",X"BD",X"DB",X"BC",X"23",X"C9",X"C0",X"BA",X"17",X"C2",X"29",X"C2",X"FF",
		X"C1",X"53",X"C2",X"1B",X"C3",X"F7",X"C2",X"02",X"00",X"01",X"C3",X"11",X"C3",X"29",X"C3",X"29",
		X"C2",X"1B",X"C3",X"F7",X"C2",X"01",X"C3",X"29",X"C3",X"29",X"C2",X"1B",X"C3",X"6F",X"C2",X"89",
		X"C3",X"7D",X"C2",X"97",X"C2",X"AF",X"C2",X"BD",X"C2",X"CF",X"C2",X"D9",X"C2",X"F7",X"C2",X"03",
		X"00",X"01",X"C3",X"29",X"C3",X"29",X"C2",X"3D",X"C2",X"0D",X"C2",X"05",X"00",X"00",X"00",X"67",
		X"BF",X"E3",X"C9",X"06",X"00",X"B3",X"C3",X"0F",X"00",X"00",X"00",X"23",X"CA",X"06",X"00",X"B3",
		X"C3",X"0F",X"00",X"00",X"00",X"63",X"CA",X"06",X"00",X"B3",X"C3",X"0F",X"00",X"00",X"00",X"A3",
		X"CA",X"05",X"00",X"B7",X"C3",X"0D",X"01",X"EB",X"C3",X"EF",X"C3",X"00",X"00",X"F1",X"CA",X"04",
		X"00",X"EF",X"C3",X"F3",X"C3",X"F3",X"C3",X"07",X"01",X"0F",X"C4",X"05",X"01",X"00",X"00",X"4F",
		X"CB",X"04",X"00",X"27",X"C4",X"0F",X"00",X"00",X"00",X"AF",X"CB",X"04",X"00",X"27",X"C4",X"0F");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
