library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_sp_bits_4 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_sp_bits_4 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"96",X"00",X"00",X"00",X"31",X"00",
		X"00",X"00",X"39",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"BA",X"AA",X"A0",X"0B",X"EB",X"AA",X"AA",X"BB",X"BB",X"AA",X"EA",
		X"BB",X"9B",X"AA",X"BE",X"BB",X"9B",X"99",X"EB",X"BA",X"BB",X"BB",X"BE",X"AA",X"B5",X"5B",X"BB",
		X"AA",X"55",X"55",X"BB",X"AA",X"55",X"55",X"B5",X"AA",X"5F",X"55",X"55",X"55",X"FF",X"FF",X"F5",
		X"AA",X"5F",X"55",X"55",X"AA",X"55",X"55",X"B5",X"AA",X"55",X"55",X"BB",X"AF",X"B5",X"5B",X"BB",
		X"BA",X"BB",X"BB",X"BE",X"BB",X"9B",X"99",X"EB",X"BB",X"9B",X"AA",X"BE",X"BB",X"BB",X"AA",X"EA",
		X"0B",X"EB",X"AA",X"AA",X"00",X"BA",X"AA",X"A0",X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"AE",X"00",X"00",
		X"BE",X"EA",X"00",X"00",X"55",X"BB",X"EA",X"00",X"55",X"55",X"5B",X"A0",X"FF",X"FF",X"FF",X"5A",
		X"55",X"55",X"5B",X"A0",X"55",X"BB",X"EA",X"00",X"BE",X"EA",X"00",X"00",X"AA",X"AE",X"00",X"00",
		X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"9B",X"AA",X"09",X"00",X"BB",X"BB",X"99",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"9B",X"00",X"00",X"BA",X"99",X"00",X"00",X"BA",X"99",X"90",X"90",X"B5",X"99",X"99",X"99",
		X"AA",X"BB",X"AA",X"90",X"AA",X"BB",X"AA",X"00",X"AA",X"55",X"AA",X"00",X"AA",X"55",X"99",X"00",
		X"AA",X"FF",X"B9",X"A0",X"AF",X"FF",X"BB",X"AA",X"BA",X"5F",X"BB",X"BA",X"BA",X"56",X"55",X"EE",
		X"BB",X"B5",X"55",X"BE",X"BB",X"BB",X"F5",X"EB",X"AB",X"AB",X"FF",X"BE",X"0A",X"AA",X"5F",X"BB",
		X"00",X"AA",X"55",X"BB",X"00",X"AA",X"B5",X"5B",X"00",X"AA",X"BB",X"F5",X"00",X"99",X"BB",X"FF",
		X"00",X"99",X"CB",X"FF",X"00",X"00",X"BE",X"5F",X"00",X"00",X"EB",X"55",X"00",X"90",X"AE",X"B5",
		X"00",X"99",X"AA",X"BB",X"00",X"09",X"AA",X"AB",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",
		X"5B",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",
		X"B5",X"A0",X"00",X"00",X"AB",X"BA",X"00",X"00",X"AA",X"BB",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"A0",X"00",X"00",X"5A",X"BA",X"00",X"00",X"55",X"BB",X"00",X"00",X"55",X"BB",X"00",X"00",
		X"A5",X"BB",X"90",X"00",X"A5",X"9B",X"90",X"00",X"A5",X"9B",X"99",X"00",X"A9",X"9B",X"09",X"00",
		X"A9",X"BB",X"09",X"00",X"A9",X"B9",X"00",X"00",X"9B",X"B9",X"00",X"00",X"9B",X"B9",X"00",X"00",
		X"9B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"5B",X"99",X"00",X"BB",X"5B",X"99",X"00",
		X"BB",X"5B",X"90",X"00",X"B9",X"55",X"A0",X"00",X"A9",X"F5",X"A9",X"00",X"AA",X"F5",X"A9",X"00",
		X"AA",X"FF",X"A9",X"00",X"AA",X"FF",X"A9",X"00",X"99",X"5F",X"AA",X"00",X"99",X"55",X"AA",X"00",
		X"99",X"B5",X"BA",X"00",X"09",X"B5",X"EA",X"00",X"09",X"BB",X"BA",X"00",X"00",X"EB",X"CA",X"00",
		X"09",X"BE",X"BA",X"00",X"09",X"EB",X"CA",X"00",X"99",X"EE",X"BA",X"00",X"99",X"AA",X"BA",X"00",
		X"99",X"AA",X"BC",X"00",X"99",X"0A",X"BB",X"00",X"09",X"0A",X"BB",X"00",X"00",X"00",X"5B",X"00",
		X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"B5",X"00",
		X"00",X"00",X"B5",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"0B",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"BB",X"BE",X"00",X"00",X"AA",X"BB",X"00",X"00",X"AA",X"BB",X"00",X"00",X"AA",X"BB",X"00",
		X"00",X"AA",X"BB",X"00",X"00",X"AA",X"AB",X"00",X"00",X"AA",X"AB",X"00",X"00",X"99",X"AB",X"00",
		X"00",X"BB",X"9B",X"00",X"00",X"B5",X"9B",X"00",X"00",X"55",X"9B",X"00",X"00",X"5F",X"BB",X"00",
		X"99",X"55",X"BB",X"00",X"99",X"5F",X"99",X"00",X"00",X"5F",X"99",X"00",X"00",X"5A",X"99",X"00",
		X"00",X"5F",X"9A",X"00",X"00",X"5F",X"9A",X"00",X"00",X"55",X"9A",X"00",X"00",X"5F",X"9A",X"00",
		X"00",X"55",X"9A",X"00",X"09",X"5F",X"99",X"00",X"99",X"55",X"9B",X"00",X"90",X"55",X"EE",X"00",
		X"00",X"55",X"EB",X"00",X"00",X"55",X"BE",X"00",X"00",X"B5",X"EB",X"00",X"00",X"55",X"BE",X"00",
		X"00",X"B5",X"EA",X"00",X"00",X"B5",X"BA",X"00",X"00",X"B5",X"A0",X"00",X"00",X"B5",X"A0",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B5",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"EB",X"00",X"00",X"00",X"E5",X"00",X"00",
		X"00",X"EB",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"AB",X"00",X"00",
		X"00",X"A5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"A5",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"05",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"05",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",
		X"00",X"50",X"00",X"30",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"3F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",
		X"05",X"00",X"00",X"FF",X"05",X"00",X"00",X"00",X"0F",X"00",X"00",X"05",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"50",X"00",X"00",X"FF",X"F0",X"00",X"00",X"F0",X"F0",X"00",X"00",X"30",
		X"F0",X"00",X"00",X"55",X"F3",X"00",X"00",X"3F",X"33",X"00",X"00",X"FF",X"3F",X"00",X"00",X"05",
		X"0F",X"35",X"50",X"0F",X"0F",X"00",X"F0",X"F0",X"0F",X"0F",X"F3",X"00",X"0F",X"0F",X"F0",X"5A",
		X"00",X"00",X"00",X"55",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"50",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"FF",X"50",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"3F",X"05",X"00",X"00",X"03",X"00",X"00",X"00",X"FF",X"30",X"00",
		X"05",X"05",X"30",X"00",X"0F",X"50",X"03",X"00",X"FF",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",
		X"F0",X"00",X"F0",X"00",X"50",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"50",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"50",X"00",X"F9",X"00",
		X"53",X"00",X"5F",X"00",X"53",X"00",X"05",X"00",X"55",X"00",X"09",X"00",X"59",X"00",X"99",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"44",X"44",X"00",X"06",X"66",X"67",X"00",X"FF",X"6F",X"66",
		X"00",X"00",X"44",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"94",X"00",X"00",X"00",
		X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"4F",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"46",X"00",X"00",X"00",
		X"4F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",
		X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"94",X"00",X"00",X"00",
		X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"5A",X"00",X"00",
		X"00",X"5A",X"00",X"00",X"00",X"A0",X"05",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"FF",X"A0",X"00",X"00",X"FF",X"E0",X"00",X"00",X"F5",X"A0",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"A0",X"55",X"00",X"00",X"5A",X"55",X"00",X"00",
		X"5A",X"55",X"00",X"00",X"F5",X"F5",X"00",X"00",X"F5",X"55",X"00",X"00",X"0F",X"F5",X"E0",X"00",
		X"00",X"5F",X"E0",X"00",X"00",X"EF",X"A0",X"00",X"00",X"E5",X"A0",X"00",X"00",X"55",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"0D",X"D9",X"00",X"00",X"00",X"9D",X"00",X"00",
		X"00",X"9D",X"90",X"00",X"09",X"99",X"90",X"00",X"E0",X"99",X"90",X"00",X"90",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"00",X"99",X"99",X"00",X"90",X"99",X"99",X"00",X"00",X"D9",X"99",X"00",
		X"00",X"D9",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",
		X"00",X"99",X"90",X"00",X"09",X"99",X"99",X"00",X"09",X"99",X"9D",X"00",X"09",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"90",X"99",X"99",X"09",
		X"99",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"90",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"E3",X"00",X"00",X"05",X"33",X"00",
		X"00",X"55",X"EE",X"00",X"00",X"5E",X"5E",X"00",X"00",X"55",X"55",X"00",X"00",X"F5",X"53",X"00",
		X"00",X"55",X"50",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"30",X"00",
		X"35",X"0F",X"30",X"00",X"55",X"50",X"30",X"00",X"F5",X"55",X"33",X"00",X"FE",X"55",X"5E",X"00",
		X"0F",X"03",X"5E",X"00",X"30",X"F3",X"55",X"00",X"55",X"EE",X"55",X"00",X"00",X"5E",X"55",X"00",
		X"0F",X"55",X"E5",X"00",X"5F",X"55",X"5E",X"00",X"00",X"03",X"55",X"00",X"00",X"F5",X"55",X"00",
		X"00",X"F5",X"55",X"00",X"00",X"5F",X"53",X"00",X"00",X"5E",X"05",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"30",X"05",X"00",X"00",X"E0",X"55",X"00",X"00",X"E3",X"55",X"00",X"00",X"5E",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"5E",X"FF",X"00",X"05",X"E5",X"FE",X"00",X"05",X"E5",X"E5",X"00",
		X"0F",X"EE",X"55",X"00",X"00",X"5F",X"55",X"00",X"00",X"F5",X"55",X"00",X"00",X"F5",X"55",X"00",
		X"00",X"55",X"F5",X"00",X"00",X"55",X"F5",X"00",X"00",X"5F",X"55",X"30",X"00",X"55",X"5E",X"30",
		X"00",X"F5",X"5E",X"30",X"00",X"5F",X"E5",X"00",X"0E",X"F5",X"5E",X"00",X"5E",X"FF",X"5E",X"00",
		X"5E",X"FF",X"5E",X"00",X"55",X"55",X"5E",X"00",X"F5",X"55",X"55",X"00",X"F5",X"F5",X"55",X"00",
		X"0F",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"F5",X"F5",X"00",
		X"00",X"E5",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"00",X"00",X"00",
		X"EB",X"99",X"00",X"00",X"E4",X"99",X"00",X"00",X"F7",X"55",X"00",X"00",X"F3",X"EE",X"99",X"00",
		X"53",X"BB",X"90",X"00",X"55",X"24",X"99",X"90",X"F5",X"77",X"E9",X"99",X"9F",X"59",X"BE",X"99",
		X"5E",X"53",X"9B",X"FF",X"59",X"39",X"99",X"EE",X"59",X"99",X"99",X"BB",X"9F",X"93",X"5F",X"FE",
		X"9F",X"33",X"FF",X"9B",X"FF",X"33",X"FF",X"B5",X"FF",X"39",X"FF",X"5F",X"FF",X"39",X"FF",X"95",
		X"F5",X"39",X"FF",X"99",X"55",X"39",X"FF",X"99",X"55",X"9F",X"FF",X"99",X"77",X"9F",X"FF",X"99",
		X"44",X"35",X"FF",X"99",X"BB",X"59",X"FF",X"99",X"FF",X"F5",X"FF",X"99",X"FF",X"99",X"5F",X"99",
		X"00",X"B9",X"95",X"95",X"00",X"BB",X"99",X"55",X"00",X"FF",X"99",X"55",X"00",X"00",X"51",X"5F",
		X"00",X"00",X"BB",X"FF",X"00",X"00",X"FF",X"44",X"00",X"00",X"5F",X"BB",X"00",X"00",X"00",X"BF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"2A",X"00",X"00",X"00",X"02",X"00",X"00",
		X"04",X"EE",X"00",X"00",X"44",X"4E",X"00",X"00",X"55",X"7E",X"00",X"00",X"35",X"74",X"00",X"00",
		X"35",X"54",X"00",X"00",X"59",X"57",X"00",X"00",X"9F",X"57",X"00",X"00",X"FF",X"F5",X"00",X"00",
		X"F5",X"F5",X"90",X"00",X"5F",X"F5",X"00",X"00",X"5F",X"55",X"90",X"00",X"5F",X"55",X"99",X"00",
		X"5F",X"55",X"90",X"00",X"55",X"55",X"99",X"00",X"75",X"99",X"90",X"00",X"75",X"99",X"99",X"00",
		X"75",X"99",X"A9",X"00",X"75",X"99",X"A9",X"00",X"47",X"99",X"A9",X"00",X"47",X"95",X"AA",X"00",
		X"E4",X"FF",X"EA",X"00",X"E4",X"FF",X"EA",X"00",X"E5",X"FF",X"EA",X"00",X"EE",X"FF",X"EA",X"00",
		X"EE",X"FF",X"EE",X"00",X"AE",X"FF",X"9E",X"00",X"AE",X"FF",X"5E",X"00",X"0A",X"FF",X"5E",X"00",
		X"0A",X"FF",X"9E",X"00",X"0A",X"FF",X"59",X"00",X"0A",X"FF",X"59",X"00",X"00",X"5F",X"55",X"00",
		X"00",X"F9",X"93",X"00",X"00",X"99",X"95",X"90",X"00",X"99",X"99",X"00",X"00",X"99",X"95",X"90",
		X"00",X"99",X"95",X"90",X"00",X"99",X"35",X"99",X"00",X"59",X"55",X"90",X"00",X"59",X"55",X"90",
		X"00",X"95",X"55",X"00",X"00",X"95",X"5E",X"90",X"00",X"E4",X"5E",X"00",X"00",X"E4",X"EA",X"90",
		X"00",X"E4",X"AA",X"00",X"00",X"04",X"55",X"00",X"00",X"AA",X"55",X"00",X"00",X"00",X"59",X"00",
		X"00",X"00",X"59",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",
		X"00",X"50",X"0F",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"B5",X"F5",X"00",
		X"00",X"55",X"F5",X"00",X"00",X"5B",X"0F",X"00",X"00",X"B5",X"55",X"00",X"00",X"BB",X"B5",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"55",X"55",X"00",X"00",X"5B",X"F0",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"5B",X"5B",X"00",X"0F",X"55",X"55",X"00",X"0F",X"BB",X"55",X"00",
		X"F5",X"55",X"B5",X"00",X"F5",X"FF",X"E5",X"00",X"BB",X"FB",X"B5",X"00",X"B5",X"B5",X"B5",X"00",
		X"BB",X"BB",X"50",X"00",X"BB",X"BB",X"00",X"00",X"B5",X"55",X"00",X"00",X"B5",X"55",X"00",X"00",
		X"F5",X"55",X"00",X"00",X"F0",X"5B",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"F5",X"B0",X"00",
		X"00",X"5F",X"5B",X"00",X"00",X"B5",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"55",X"B0",X"00",X"BB",X"5F",X"B0",X"00",X"BB",X"BB",X"B0",X"00",X"55",X"55",X"00",X"00",
		X"BB",X"55",X"00",X"00",X"5B",X"B5",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"55",X"00",X"00",
		X"B0",X"B5",X"00",X"00",X"B0",X"BB",X"00",X"00",X"B0",X"5F",X"00",X"00",X"B0",X"5F",X"00",X"00",
		X"B0",X"5F",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"90",X"00",
		X"99",X"99",X"59",X"00",X"9A",X"A9",X"95",X"00",X"93",X"A9",X"99",X"90",X"A4",X"99",X"AA",X"90",
		X"77",X"99",X"FA",X"44",X"75",X"59",X"9A",X"A3",X"55",X"55",X"FA",X"AA",X"F3",X"55",X"F9",X"5A",
		X"53",X"F5",X"99",X"4A",X"35",X"F5",X"F9",X"5A",X"35",X"95",X"F9",X"9A",X"35",X"F5",X"F9",X"99",
		X"33",X"F5",X"59",X"99",X"33",X"5F",X"59",X"9A",X"53",X"FF",X"59",X"5A",X"55",X"FF",X"99",X"5A",
		X"75",X"FF",X"F9",X"A5",X"45",X"55",X"FF",X"A5",X"47",X"59",X"99",X"A3",X"47",X"99",X"FF",X"44",
		X"44",X"99",X"51",X"EA",X"EE",X"A0",X"AE",X"AA",X"99",X"99",X"AA",X"00",X"39",X"FF",X"95",X"00",
		X"00",X"F9",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"09",X"09",X"99",X"09",X"99",X"99",X"90",
		X"55",X"99",X"99",X"59",X"EE",X"EE",X"EE",X"EE",X"BB",X"BB",X"BB",X"BB",X"44",X"5F",X"99",X"55",
		X"77",X"95",X"9F",X"FE",X"45",X"99",X"FF",X"5B",X"55",X"99",X"FF",X"B5",X"FF",X"99",X"FF",X"9B",
		X"E5",X"99",X"FF",X"99",X"EE",X"39",X"FF",X"99",X"F5",X"39",X"FF",X"99",X"F5",X"39",X"FF",X"99",
		X"F5",X"39",X"FF",X"99",X"FF",X"39",X"FF",X"99",X"FF",X"39",X"FF",X"99",X"FF",X"39",X"FF",X"99",
		X"F5",X"39",X"FF",X"9E",X"55",X"33",X"FF",X"55",X"55",X"93",X"FF",X"55",X"77",X"95",X"9F",X"55",
		X"44",X"5F",X"99",X"55",X"BF",X"BB",X"BB",X"BB",X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"F9",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"C9",X"99",X"99",X"00",
		X"BC",X"9C",X"99",X"00",X"B6",X"C0",X"CC",X"90",X"AA",X"BE",X"BE",X"90",X"AC",X"9B",X"90",X"99",
		X"AA",X"9B",X"EC",X"94",X"BE",X"9B",X"BE",X"F4",X"EB",X"95",X"EB",X"54",X"BE",X"9B",X"BB",X"59",
		X"BB",X"95",X"BB",X"59",X"EE",X"9B",X"BB",X"59",X"5F",X"9F",X"BB",X"59",X"BB",X"9B",X"BB",X"59",
		X"BB",X"9F",X"BB",X"59",X"BB",X"9F",X"BB",X"59",X"6F",X"9F",X"FB",X"54",X"B6",X"9F",X"BF",X"F4",
		X"9B",X"9B",X"F9",X"94",X"C9",X"BB",X"BB",X"90",X"BB",X"BB",X"BB",X"90",X"B6",X"C0",X"CC",X"00",
		X"BC",X"9C",X"99",X"00",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"E9",X"99",X"99",X"00",X"E9",X"09",X"59",X"00",X"17",X"99",X"59",X"90",
		X"17",X"99",X"22",X"99",X"19",X"A9",X"D2",X"99",X"99",X"77",X"9E",X"00",X"50",X"D7",X"A9",X"00",
		X"9E",X"7D",X"A9",X"99",X"E9",X"77",X"A9",X"FE",X"E9",X"77",X"A9",X"99",X"5E",X"77",X"AE",X"FE",
		X"59",X"77",X"AE",X"00",X"99",X"77",X"EE",X"00",X"19",X"70",X"D2",X"00",X"17",X"00",X"22",X"00",
		X"16",X"00",X"50",X"00",X"E9",X"00",X"50",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A9",X"AA",X"AA",X"AA",
		X"99",X"7A",X"99",X"99",X"9A",X"EA",X"99",X"99",X"A3",X"AE",X"99",X"FF",X"A3",X"EA",X"93",X"99",
		X"3A",X"99",X"33",X"99",X"A3",X"93",X"7A",X"99",X"99",X"39",X"AA",X"9E",X"FF",X"9F",X"A9",X"9E",
		X"F9",X"FA",X"99",X"9E",X"FF",X"FA",X"99",X"9E",X"F9",X"99",X"99",X"95",X"FF",X"95",X"53",X"9E",
		X"F9",X"99",X"AA",X"9E",X"FF",X"F9",X"AA",X"95",X"F9",X"F9",X"AA",X"EE",X"FF",X"EF",X"AA",X"95",
		X"99",X"EE",X"EA",X"95",X"3A",X"9E",X"5A",X"9E",X"A3",X"99",X"EA",X"99",X"3A",X"EE",X"9E",X"99",
		X"3E",X"EA",X"99",X"99",X"9E",X"AE",X"99",X"FF",X"99",X"EA",X"99",X"99",X"D9",X"5A",X"99",X"99",
		X"0D",X"D9",X"D9",X"D9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"3E",X"99",X"00",
		X"99",X"EE",X"99",X"00",X"99",X"99",X"99",X"00",X"FF",X"FF",X"99",X"00",X"99",X"99",X"AA",X"00",
		X"A7",X"A7",X"AA",X"00",X"AA",X"AA",X"A9",X"00",X"AA",X"AA",X"95",X"00",X"AA",X"AA",X"99",X"00",
		X"A9",X"AA",X"99",X"00",X"A4",X"AA",X"99",X"00",X"AA",X"AA",X"99",X"00",X"AA",X"AA",X"99",X"00",
		X"AA",X"AA",X"99",X"00",X"AA",X"AA",X"99",X"00",X"A9",X"AA",X"99",X"00",X"A4",X"AA",X"99",X"00",
		X"EA",X"AA",X"99",X"00",X"AE",X"AA",X"05",X"00",X"EE",X"AE",X"A0",X"00",X"EE",X"E5",X"AA",X"00",
		X"99",X"99",X"AA",X"00",X"FF",X"FF",X"99",X"00",X"99",X"99",X"99",X"00",X"D9",X"EE",X"99",X"00",
		X"00",X"3E",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"A9",
		X"9E",X"AA",X"AA",X"A3",X"9E",X"AA",X"EE",X"99",X"95",X"99",X"55",X"55",X"9E",X"99",X"50",X"99",
		X"99",X"99",X"99",X"39",X"99",X"49",X"33",X"A3",X"99",X"99",X"EB",X"E9",X"44",X"93",X"3E",X"99",
		X"99",X"93",X"EE",X"09",X"AA",X"90",X"3E",X"A9",X"AA",X"90",X"EB",X"E9",X"AA",X"00",X"EA",X"A9",
		X"AA",X"93",X"EB",X"E9",X"44",X"A3",X"EE",X"99",X"EE",X"99",X"EB",X"39",X"9E",X"49",X"3B",X"A3",
		X"99",X"E9",X"99",X"39",X"99",X"99",X"55",X"99",X"9E",X"99",X"55",X"55",X"9E",X"AA",X"EE",X"9E",
		X"9E",X"AA",X"EA",X"99",X"99",X"99",X"99",X"E9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",
		X"E3",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"EA",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"39",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"90",X"90",X"99",X"99",X"09",X"09",X"22",X"29",X"99",X"99",X"22",X"22",
		X"99",X"99",X"22",X"22",X"33",X"A9",X"22",X"22",X"13",X"39",X"22",X"22",X"A1",X"A9",X"22",X"22",
		X"1A",X"F9",X"22",X"22",X"92",X"22",X"22",X"22",X"23",X"77",X"22",X"22",X"71",X"47",X"22",X"22",
		X"13",X"47",X"22",X"22",X"19",X"44",X"22",X"22",X"19",X"44",X"22",X"22",X"19",X"44",X"22",X"22",
		X"99",X"44",X"22",X"22",X"72",X"44",X"22",X"22",X"11",X"77",X"22",X"22",X"12",X"47",X"22",X"22",
		X"11",X"77",X"22",X"22",X"77",X"47",X"22",X"22",X"23",X"77",X"22",X"22",X"92",X"22",X"22",X"22",
		X"1A",X"F9",X"22",X"22",X"A1",X"29",X"22",X"22",X"13",X"29",X"22",X"22",X"3A",X"A9",X"22",X"22",
		X"99",X"00",X"22",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"33",X"00",X"00",
		X"90",X"39",X"00",X"00",X"90",X"39",X"00",X"00",X"90",X"39",X"00",X"00",X"90",X"39",X"00",X"00",
		X"90",X"39",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"33",X"33",X"00",X"00",X"90",X"39",X"00",X"00",
		X"90",X"39",X"00",X"00",X"90",X"39",X"00",X"00",X"90",X"39",X"00",X"00",X"90",X"39",X"00",X"00",
		X"99",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"09",X"00",X"90",X"99",
		X"99",X"09",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"DD",X"22",X"22",X"11",
		X"11",X"99",X"91",X"11",X"11",X"19",X"31",X"11",X"F7",X"91",X"11",X"99",X"11",X"91",X"77",X"99",
		X"11",X"31",X"77",X"99",X"ED",X"31",X"77",X"99",X"44",X"31",X"77",X"99",X"44",X"31",X"77",X"99",
		X"44",X"31",X"77",X"99",X"44",X"31",X"77",X"99",X"54",X"31",X"77",X"99",X"7F",X"31",X"77",X"95",
		X"1D",X"91",X"77",X"59",X"EE",X"91",X"57",X"99",X"11",X"91",X"11",X"99",X"11",X"19",X"30",X"11",
		X"77",X"99",X"91",X"11",X"52",X"20",X"22",X"11",X"22",X"22",X"25",X"22",X"99",X"00",X"22",X"22",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"09",X"00",
		X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"90",
		X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"99",X"99",X"90",
		X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"09",X"00",X"09",X"99",X"00",X"00",
		X"30",X"30",X"05",X"00",X"30",X"E0",X"55",X"55",X"53",X"E3",X"55",X"55",X"53",X"5E",X"55",X"55",
		X"55",X"55",X"55",X"55",X"55",X"5E",X"FF",X"55",X"55",X"E5",X"FE",X"55",X"55",X"E5",X"E5",X"55",
		X"5F",X"5E",X"55",X"55",X"55",X"5F",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"F5",X"55",X"55",
		X"55",X"55",X"F5",X"55",X"55",X"55",X"F5",X"55",X"55",X"5F",X"55",X"55",X"55",X"55",X"5E",X"55",
		X"55",X"F5",X"5E",X"55",X"55",X"5F",X"E5",X"55",X"5F",X"F5",X"5E",X"55",X"5E",X"FF",X"5E",X"55",
		X"5E",X"5F",X"55",X"55",X"55",X"55",X"5E",X"55",X"F5",X"55",X"55",X"55",X"F5",X"F5",X"55",X"55",
		X"5F",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"F5",X"55",
		X"55",X"E5",X"55",X"55",X"53",X"E5",X"55",X"55",X"30",X"E3",X"55",X"55",X"00",X"00",X"53",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",
		X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",
		X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",
		X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"09",X"00",X"00",
		X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",
		X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",
		X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",
		X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"19",X"11",X"00",X"00",X"01",X"11",X"00",X"00",
		X"01",X"11",X"10",X"00",X"01",X"11",X"90",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"F0",X"00",X"00",X"11",X"0F",X"11",X"00",X"11",X"60",X"00",X"00",
		X"11",X"66",X"00",X"00",X"00",X"D9",X"02",X"00",X"02",X"19",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"19",X"90",X"00",X"00",X"10",X"19",X"00",X"00",X"10",X"19",X"00",X"00",X"10",X"11",X"00",
		X"00",X"10",X"01",X"00",X"01",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"99",X"19",X"00",X"00",X"99",X"10",X"09",X"00",X"00",X"00",X"11",X"00",X"00",X"F0",X"11",X"00",
		X"09",X"99",X"19",X"00",X"99",X"F9",X"F1",X"00",X"99",X"66",X"D1",X"10",X"11",X"FF",X"D1",X"10",
		X"11",X"F6",X"D1",X"90",X"00",X"00",X"D0",X"00",X"11",X"00",X"01",X"00",X"11",X"0D",X"19",X"00",
		X"19",X"91",X"10",X"00",X"09",X"91",X"11",X"00",X"00",X"91",X"11",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"00",X"00",X"00",X"09",X"20",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"01",X"00",X"00",X"11",X"00",X"01",X"11",X"11",X"00",
		X"00",X"00",X"10",X"00",X"00",X"01",X"00",X"06",X"01",X"01",X"00",X"00",X"00",X"11",X"0F",X"60",
		X"00",X"00",X"FF",X"99",X"00",X"60",X"09",X"99",X"44",X"06",X"00",X"FF",X"44",X"00",X"00",X"0F",
		X"11",X"11",X"60",X"0F",X"94",X"66",X"00",X"6F",X"09",X"66",X"66",X"F0",X"00",X"10",X"06",X"00",
		X"00",X"10",X"66",X"00",X"00",X"06",X"00",X"00",X"04",X"66",X"00",X"05",X"41",X"44",X"00",X"50",
		X"44",X"11",X"00",X"90",X"40",X"14",X"00",X"55",X"09",X"11",X"01",X"94",X"90",X"10",X"90",X"19",
		X"00",X"90",X"11",X"19",X"00",X"90",X"44",X"14",X"00",X"90",X"99",X"14",X"00",X"00",X"90",X"01",
		X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",
		X"00",X"44",X"40",X"00",X"00",X"40",X"40",X"00",X"40",X"00",X"40",X"00",X"44",X"00",X"40",X"00",
		X"44",X"00",X"40",X"00",X"44",X"00",X"00",X"00",X"04",X"40",X"00",X"00",X"11",X"40",X"00",X"00",
		X"01",X"04",X"00",X"00",X"11",X"04",X"00",X"00",X"00",X"11",X"09",X"00",X"60",X"11",X"10",X"00",
		X"60",X"00",X"14",X"00",X"50",X"00",X"11",X"00",X"65",X"06",X"14",X"00",X"65",X"66",X"10",X"00",
		X"60",X"00",X"00",X"00",X"69",X"66",X"99",X"00",X"99",X"00",X"44",X"00",X"00",X"00",X"11",X"00",
		X"06",X"66",X"11",X"00",X"00",X"00",X"44",X"44",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"11",X"91",X"00",
		X"00",X"01",X"09",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"63",X"00",X"00",X"00",X"64",X"00",X"00",
		X"00",X"33",X"00",X"00",X"30",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"03",X"31",X"00",X"00",
		X"03",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"41",X"03",X"00",X"03",X"46",X"33",X"00",
		X"00",X"F6",X"39",X"00",X"00",X"FF",X"33",X"00",X"00",X"FF",X"09",X"00",X"30",X"4F",X"00",X"00",
		X"03",X"FF",X"00",X"00",X"33",X"F6",X"39",X"00",X"03",X"66",X"30",X"00",X"36",X"66",X"13",X"00",
		X"33",X"16",X"33",X"00",X"30",X"36",X"33",X"00",X"30",X"33",X"39",X"00",X"00",X"33",X"39",X"00",
		X"03",X"30",X"03",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"90",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"00",X"11",X"99",X"99",X"99",X"16",X"99",X"99",X"39",X"66",X"99",X"09",
		X"31",X"F6",X"36",X"00",X"61",X"61",X"66",X"00",X"66",X"16",X"31",X"00",X"3F",X"41",X"61",X"00",
		X"61",X"FF",X"11",X"00",X"96",X"FF",X"99",X"00",X"36",X"F4",X"99",X"00",X"66",X"FF",X"99",X"00",
		X"64",X"4F",X"99",X"00",X"66",X"46",X"99",X"00",X"66",X"41",X"19",X"00",X"91",X"61",X"19",X"00",
		X"99",X"61",X"66",X"00",X"66",X"66",X"63",X"00",X"16",X"66",X"99",X"00",X"63",X"96",X"99",X"00",
		X"66",X"99",X"99",X"90",X"69",X"09",X"99",X"90",X"00",X"30",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"39",X"99",X"00",X"00",X"33",X"69",X"00",
		X"99",X"93",X"61",X"00",X"00",X"93",X"13",X"00",X"99",X"99",X"39",X"00",X"00",X"91",X"33",X"00",
		X"03",X"91",X"33",X"00",X"03",X"16",X"93",X"39",X"99",X"66",X"13",X"39",X"99",X"66",X"39",X"30",
		X"19",X"69",X"39",X"00",X"11",X"11",X"99",X"00",X"63",X"63",X"91",X"00",X"33",X"16",X"99",X"00",
		X"13",X"66",X"99",X"30",X"03",X"91",X"93",X"30",X"33",X"44",X"39",X"00",X"34",X"66",X"19",X"00",
		X"33",X"61",X"11",X"00",X"33",X"61",X"39",X"00",X"63",X"11",X"99",X"00",X"10",X"19",X"93",X"00",
		X"93",X"99",X"19",X"00",X"00",X"69",X"61",X"00",X"03",X"39",X"66",X"30",X"33",X"63",X"91",X"30",
		X"36",X"99",X"99",X"00",X"90",X"99",X"33",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"90",X"96",X"09",X"00",
		X"90",X"36",X"93",X"00",X"09",X"61",X"30",X"00",X"99",X"13",X"00",X"00",X"99",X"33",X"93",X"00",
		X"99",X"99",X"33",X"00",X"11",X"96",X"33",X"00",X"06",X"11",X"63",X"00",X"33",X"13",X"13",X"00",
		X"33",X"93",X"99",X"90",X"01",X"13",X"99",X"00",X"16",X"39",X"93",X"00",X"41",X"69",X"33",X"00",
		X"90",X"99",X"99",X"00",X"69",X"33",X"39",X"00",X"34",X"63",X"33",X"00",X"30",X"11",X"33",X"00",
		X"46",X"31",X"93",X"00",X"46",X"33",X"99",X"00",X"91",X"99",X"99",X"00",X"31",X"39",X"33",X"00",
		X"99",X"31",X"33",X"00",X"36",X"36",X"33",X"90",X"03",X"10",X"93",X"90",X"00",X"99",X"93",X"90",
		X"99",X"99",X"93",X"00",X"09",X"33",X"99",X"00",X"30",X"09",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"00",X"00",X"33",X"00",X"00",X"90",X"30",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"39",X"00",X"00",X"03",X"39",X"00",X"00",X"33",X"39",X"00",X"00",X"00",X"33",X"00",X"90",
		X"00",X"93",X"99",X"00",X"03",X"99",X"33",X"30",X"33",X"93",X"33",X"30",X"33",X"93",X"33",X"00",
		X"33",X"33",X"33",X"00",X"33",X"33",X"99",X"00",X"39",X"33",X"33",X"00",X"09",X"33",X"99",X"00",
		X"03",X"33",X"90",X"00",X"33",X"33",X"30",X"00",X"99",X"33",X"00",X"00",X"99",X"33",X"90",X"00",
		X"09",X"33",X"93",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"33",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"03",X"90",X"00",
		X"55",X"00",X"30",X"00",X"55",X"33",X"30",X"00",X"05",X"03",X"03",X"00",X"35",X"03",X"39",X"00",
		X"35",X"03",X"39",X"00",X"33",X"F3",X"39",X"00",X"00",X"33",X"93",X"00",X"05",X"39",X"33",X"90",
		X"55",X"99",X"33",X"00",X"55",X"99",X"53",X"00",X"55",X"99",X"35",X"00",X"53",X"99",X"39",X"00",
		X"39",X"99",X"53",X"00",X"03",X"99",X"03",X"00",X"33",X"99",X"03",X"00",X"59",X"99",X"53",X"00",
		X"50",X"99",X"33",X"00",X"00",X"39",X"30",X"00",X"00",X"03",X"90",X"00",X"05",X"09",X"90",X"00",
		X"05",X"90",X"39",X"00",X"50",X"00",X"39",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"60",X"00",
		X"00",X"FF",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"10",X"00",
		X"00",X"FF",X"61",X"00",X"00",X"55",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"07",X"FF",X"40",X"00",
		X"77",X"FF",X"46",X"00",X"07",X"5A",X"64",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"7F",X"55",X"00",X"00",X"77",X"FF",X"60",X"00",
		X"77",X"FF",X"61",X"00",X"7F",X"5A",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"5A",X"00",X"00",X"5F",X"55",X"00",X"00",X"5F",X"FF",X"60",X"00",
		X"5F",X"FF",X"61",X"00",X"FF",X"5A",X"16",X"22",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"5A",X"00",X"00",X"5F",X"55",X"44",X"40",X"5F",X"FF",X"60",X"00",
		X"5F",X"FF",X"44",X"00",X"FF",X"5A",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"96",X"00",X"00",
		X"00",X"69",X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"69",X"49",X"00",
		X"00",X"96",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"05",X"00",X"00",X"3F",X"FF",X"00",X"00",X"E4",X"F5",X"00",
		X"00",X"F4",X"5F",X"00",X"00",X"F4",X"50",X"00",X"00",X"44",X"30",X"00",X"00",X"46",X"35",X"00",
		X"00",X"66",X"35",X"00",X"3F",X"6F",X"55",X"00",X"03",X"6F",X"53",X"00",X"00",X"6F",X"4F",X"00",
		X"0E",X"66",X"04",X"00",X"00",X"44",X"00",X"00",X"00",X"F4",X"00",X"00",X"00",X"44",X"F0",X"00",
		X"00",X"4F",X"F0",X"00",X"00",X"4F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"3F",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"5F",X"05",X"00",X"00",X"3F",X"FF",X"00",X"00",X"EF",X"F5",X"00",
		X"00",X"FF",X"5F",X"00",X"00",X"FF",X"50",X"00",X"00",X"FF",X"30",X"00",X"00",X"F4",X"35",X"00",
		X"00",X"F6",X"35",X"00",X"3F",X"6F",X"55",X"00",X"03",X"6F",X"53",X"00",X"00",X"4F",X"4F",X"00",
		X"0E",X"46",X"EF",X"00",X"0E",X"FF",X"FF",X"00",X"00",X"FF",X"3E",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"EF",X"F3",X"00",X"00",X"EF",X"EE",X"00",X"00",X"5F",X"00",X"00",X"00",X"3F",X"05",X"00",
		X"00",X"EE",X"05",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"5E",X"00",
		X"00",X"55",X"5E",X"00",X"00",X"55",X"F5",X"00",X"00",X"35",X"FF",X"00",X"00",X"EE",X"55",X"00",
		X"05",X"F3",X"5F",X"00",X"05",X"FF",X"55",X"00",X"05",X"53",X"35",X"00",X"35",X"53",X"35",X"00",
		X"35",X"3F",X"35",X"00",X"33",X"55",X"55",X"00",X"03",X"F3",X"53",X"00",X"00",X"F3",X"3F",X"00",
		X"0E",X"5F",X"EF",X"00",X"0E",X"F5",X"FF",X"00",X"EE",X"F5",X"3E",X"00",X"E5",X"F5",X"FE",X"00",
		X"E5",X"EF",X"53",X"00",X"00",X"EF",X"EE",X"00",X"E0",X"5F",X"F5",X"00",X"00",X"3F",X"55",X"00",
		X"E0",X"EE",X"55",X"00",X"00",X"55",X"F0",X"00",X"00",X"FF",X"F0",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"E0",X"00",X"0E",X"EE",X"E0",X"00",
		X"0E",X"33",X"EE",X"00",X"0E",X"55",X"FE",X"00",X"EE",X"FF",X"F5",X"00",X"E5",X"F3",X"F5",X"00",
		X"E5",X"55",X"F3",X"00",X"55",X"F5",X"FF",X"00",X"5E",X"55",X"5F",X"00",X"5F",X"F5",X"FF",X"00",
		X"55",X"F5",X"F5",X"00",X"55",X"FF",X"FF",X"00",X"55",X"55",X"35",X"00",X"F5",X"FF",X"5E",X"00",
		X"55",X"FF",X"33",X"00",X"53",X"F3",X"33",X"00",X"53",X"F5",X"55",X"00",X"33",X"55",X"F5",X"00",
		X"EE",X"55",X"F5",X"00",X"E5",X"FF",X"F5",X"00",X"E5",X"3F",X"F5",X"00",X"E5",X"55",X"5E",X"00",
		X"E5",X"55",X"EE",X"00",X"E5",X"E3",X"30",X"00",X"EE",X"E0",X"E0",X"00",X"0E",X"E0",X"00",X"30",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A4",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"A6",X"00",X"00",X"00",X"66",X"64",X"00",X"00",X"44",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A4",X"16",X"40",X"00",
		X"A4",X"64",X"00",X"00",X"66",X"40",X"00",X"00",X"46",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"A6",X"40",X"00",X"00",X"66",X"60",X"00",X"00",
		X"11",X"06",X"00",X"00",X"60",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"16",X"00",X"00",
		X"46",X"01",X"00",X"00",X"60",X"00",X"00",X"00",X"44",X"60",X"00",X"00",X"66",X"66",X"00",X"00",
		X"AA",X"11",X"00",X"00",X"A6",X"06",X"10",X"00",X"16",X"01",X"00",X"00",X"61",X"60",X"66",X"00",
		X"46",X"06",X"00",X"00",X"44",X"61",X"00",X"00",X"40",X"10",X"06",X"00",X"46",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"41",X"16",X"00",X"00",X"66",X"61",X"00",X"00",X"66",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"66",X"00",X"00",X"00",X"46",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"46",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"66",X"61",X"00",X"00",X"41",X"16",X"00",X"00",X"46",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"40",X"10",X"06",X"00",X"44",X"61",X"00",X"66",X"46",X"06",X"00",X"00",
		X"61",X"60",X"00",X"00",X"16",X"01",X"00",X"00",X"A6",X"06",X"10",X"00",X"AA",X"00",X"00",X"00",
		X"66",X"66",X"00",X"00",X"44",X"60",X"00",X"00",X"60",X"00",X"66",X"00",X"46",X"01",X"00",X"00",
		X"66",X"10",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"A6",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"44",X"16",X"00",X"00",
		X"44",X"01",X"00",X"00",X"46",X"00",X"00",X"00",X"66",X"40",X"00",X"00",X"A4",X"00",X"00",X"00",
		X"A4",X"16",X"40",X"00",X"66",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"44",X"46",X"00",X"00",
		X"A0",X"44",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"64",X"00",X"00",X"A6",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"A4",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"6E",X"90",X"09",X"00",X"6E",X"99",X"00",X"00",X"EE",X"90",X"90",X"00",X"E9",X"99",X"09",X"00",
		X"59",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"79",X"99",X"00",X"09",X"D7",X"99",X"00",
		X"00",X"DD",X"99",X"00",X"70",X"DD",X"D9",X"00",X"00",X"7D",X"DD",X"00",X"77",X"D7",X"DD",X"00",
		X"67",X"77",X"A2",X"00",X"07",X"77",X"99",X"00",X"06",X"DA",X"99",X"00",X"00",X"0A",X"99",X"00",
		X"00",X"0D",X"59",X"00",X"00",X"06",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"59",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DA",X"99",
		X"00",X"00",X"DA",X"99",X"00",X"00",X"A0",X"F9",X"00",X"00",X"A0",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"0D",X"AE",X"00",
		X"00",X"DD",X"AE",X"90",X"09",X"77",X"A9",X"00",X"09",X"77",X"A9",X"00",X"05",X"7D",X"DA",X"00",
		X"01",X"D7",X"DD",X"00",X"01",X"22",X"DD",X"00",X"0D",X"12",X"77",X"00",X"00",X"11",X"09",X"00",
		X"00",X"51",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"17",X"00",X"00",X"00",X"D7",X"00",X"00",
		X"09",X"D7",X"00",X"00",X"99",X"76",X"00",X"00",X"F9",X"60",X"00",X"00",X"99",X"70",X"00",X"00",
		X"00",X"99",X"99",X"99",X"0B",X"99",X"99",X"99",X"0B",X"90",X"00",X"00",X"BB",X"66",X"00",X"00",
		X"00",X"44",X"66",X"00",X"00",X"4A",X"44",X"A0",X"0B",X"EB",X"AA",X"AA",X"BB",X"55",X"AE",X"EA",
		X"BB",X"55",X"AE",X"0E",X"F4",X"55",X"11",X"00",X"F4",X"55",X"1B",X"EE",X"FF",X"55",X"11",X"EE",
		X"4F",X"55",X"11",X"EE",X"FF",X"11",X"FF",X"EE",X"11",X"FF",X"55",X"50",X"16",X"FF",X"11",X"F0",
		X"4F",X"FF",X"15",X"55",X"6F",X"F1",X"10",X"B5",X"66",X"FF",X"F0",X"BB",X"40",X"FF",X"FB",X"EE",
		X"00",X"1F",X"FF",X"EE",X"06",X"1F",X"9F",X"EE",X"60",X"11",X"AF",X"BE",X"00",X"66",X"A0",X"EA",
		X"06",X"66",X"10",X"AA",X"06",X"11",X"10",X"A0",X"BB",X"91",X"11",X"00",X"B0",X"91",X"60",X"00",
		X"00",X"91",X"00",X"00",X"00",X"90",X"00",X"60",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",
		X"00",X"06",X"00",X"06",X"00",X"00",X"00",X"66",X"00",X"00",X"10",X"66",X"00",X"00",X"11",X"66",
		X"00",X"00",X"01",X"66",X"00",X"00",X"61",X"41",X"00",X"00",X"61",X"11",X"00",X"00",X"66",X"1F",
		X"00",X"00",X"06",X"11",X"00",X"00",X"00",X"51",X"00",X"09",X"40",X"11",X"00",X"06",X"44",X"15",
		X"00",X"06",X"FF",X"16",X"00",X"10",X"FF",X"51",X"00",X"01",X"FF",X"16",X"00",X"01",X"1A",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"60",X"11",X"00",X"B0",X"60",X"10",X"00",X"00",X"60",X"00",X"00",X"00",
		X"61",X"00",X"00",X"00",X"16",X"BB",X"BB",X"00",X"66",X"BB",X"E0",X"00",X"66",X"B1",X"1E",X"00",
		X"00",X"60",X"6F",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"01",X"F0",X"66",X"00",X"11",X"66",X"F6",
		X"00",X"00",X"66",X"F6",X"00",X"00",X"66",X"F6",X"00",X"00",X"66",X"FF",X"01",X"00",X"00",X"66",
		X"00",X"00",X"00",X"66",X"00",X"01",X"66",X"66",X"00",X"00",X"61",X"16",X"00",X"00",X"01",X"11",
		X"00",X"00",X"01",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"01",X"00",X"00",X"00",X"01",
		X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"A0",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"41",X"00",X"00",X"66",X"11",X"00",X"00",X"61",X"66",X"00",X"00",X"16",X"00",X"00",X"00",
		X"66",X"11",X"11",X"E0",X"11",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"61",X"00",X"00",X"00",
		X"66",X"60",X"00",X"00",X"11",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",
		X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",
		X"00",X"00",X"00",X"61",X"00",X"00",X"11",X"61",X"00",X"00",X"11",X"61",X"00",X"00",X"11",X"11",
		X"00",X"00",X"01",X"11",X"00",X"00",X"61",X"16",X"00",X"01",X"66",X"66",X"00",X"00",X"01",X"66",
		X"01",X"00",X"01",X"66",X"00",X"00",X"66",X"FF",X"00",X"00",X"66",X"F6",X"00",X"00",X"66",X"F6",
		X"00",X"11",X"66",X"F1",X"00",X"01",X"F0",X"66",X"00",X"00",X"FF",X"FF",X"00",X"60",X"6F",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"66",X"00",X"00",X"66",X"60",X"00",X"00",
		X"61",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"11",X"11",X"E0",
		X"16",X"00",X"00",X"00",X"61",X"66",X"00",X"00",X"66",X"11",X"00",X"00",X"11",X"41",X"00",X"00",
		X"00",X"01",X"1A",X"FF",X"00",X"01",X"FF",X"16",X"00",X"10",X"FF",X"61",X"00",X"06",X"FF",X"65",
		X"00",X"06",X"44",X"65",X"00",X"09",X"40",X"65",X"00",X"00",X"00",X"65",X"00",X"00",X"06",X"66",
		X"00",X"00",X"66",X"56",X"00",X"00",X"61",X"16",X"00",X"00",X"61",X"41",X"00",X"00",X"01",X"66",
		X"06",X"00",X"11",X"66",X"00",X"00",X"10",X"66",X"00",X"00",X"00",X"66",X"00",X"06",X"00",X"06",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"66",X"B1",X"1E",X"00",X"66",X"00",X"E0",X"00",X"16",X"BB",X"00",X"00",X"61",X"00",X"00",X"00",
		X"11",X"60",X"00",X"00",X"11",X"16",X"00",X"00",X"61",X"11",X"00",X"00",X"66",X"00",X"00",X"00",
		X"11",X"00",X"60",X"00",X"44",X"11",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"10",X"03",X"00",X"00",X"10",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"10",X"06",X"00",X"00",X"10",X"06",
		X"00",X"00",X"00",X"66",X"00",X"00",X"01",X"31",X"00",X"00",X"01",X"33",X"00",X"00",X"00",X"33",
		X"00",X"00",X"06",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"40",X"03",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"3F",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"13",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"36",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"44",X"10",X"00",X"00",X"33",X"00",X"60",X"00",
		X"66",X"00",X"00",X"00",X"03",X"11",X"00",X"00",X"11",X"16",X"00",X"00",X"00",X"60",X"00",X"00",
		X"60",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"63",X"01",X"10",X"00",
		X"00",X"60",X"33",X"30",X"00",X"00",X"33",X"30",X"00",X"01",X"00",X"00",X"00",X"11",X"06",X"00",
		X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"33",X"00",X"00",X"01",X"33",
		X"00",X"00",X"00",X"33",X"00",X"01",X"66",X"33",X"00",X"00",X"61",X"06",X"00",X"00",X"01",X"00",
		X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"60",X"00",X"00",X"11",X"61",X"00",X"00",X"00",X"61",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"03",X"41",X"00",X"00",X"00",X"13",X"00",X"00",X"33",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"11",X"11",X"00",X"00",X"00",X"00",X"00",X"03",X"11",X"00",X"00",X"03",X"00",X"00",X"00",
		X"33",X"60",X"00",X"00",X"30",X"36",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"01",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"A0",X"00",X"5F",X"99",X"A0",
		X"00",X"99",X"9F",X"00",X"05",X"99",X"F9",X"BA",X"55",X"99",X"FF",X"BB",X"FF",X"99",X"FF",X"9A",
		X"55",X"99",X"FF",X"5A",X"55",X"39",X"FF",X"5A",X"53",X"39",X"FF",X"5A",X"33",X"39",X"FF",X"5A",
		X"33",X"39",X"FF",X"5A",X"53",X"39",X"FF",X"5A",X"55",X"39",X"FF",X"5A",X"55",X"39",X"FF",X"5A",
		X"FF",X"33",X"FF",X"9A",X"55",X"33",X"FF",X"5A",X"55",X"93",X"F9",X"9A",X"BB",X"99",X"9F",X"00",
		X"00",X"5F",X"99",X"0A",X"00",X"EE",X"EE",X"A0",X"B0",X"00",X"BA",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"AB",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"AB",X"00",X"00",X"00",X"B0",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"0A",X"99",X"F9",X"00",X"AA",X"99",X"FF",X"00",X"FF",X"99",X"FF",X"00",
		X"55",X"99",X"FF",X"A0",X"55",X"39",X"FF",X"A0",X"53",X"39",X"FF",X"00",X"33",X"39",X"FF",X"00",
		X"33",X"39",X"FF",X"00",X"53",X"39",X"FF",X"00",X"05",X"39",X"FF",X"50",X"05",X"39",X"FF",X"00",
		X"00",X"33",X"FF",X"00",X"00",X"33",X"FF",X"00",X"00",X"93",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"AA",X"00",X"00",X"A0",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"A0",X"BB",X"B0",X"00",X"0B",X"00",X"BB",X"00",X"00",X"AA",X"00",X"00",
		X"BB",X"99",X"00",X"00",X"05",X"39",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"39",X"F0",X"00",
		X"00",X"39",X"F0",X"00",X"53",X"39",X"F0",X"00",X"00",X"39",X"F0",X"00",X"B5",X"39",X"F0",X"B0",
		X"00",X"33",X"F0",X"B0",X"00",X"33",X"00",X"B0",X"0B",X"00",X"00",X"00",X"0B",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"B0",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"B0",X"0A",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"39",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"61",X"00",X"00",
		X"00",X"61",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"39",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"AB",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"B0",X"0B",X"00",X"BB",X"B0",X"BB",X"00",X"0B",X"B0",X"B0",X"00",X"BB",X"B0",X"B0",X"00",
		X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"BB",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"AB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"B0",X"BB",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"B0",X"00",
		X"BB",X"B0",X"B0",X"00",X"0B",X"B0",X"B0",X"00",X"BB",X"B0",X"BB",X"00",X"BB",X"B0",X"0B",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",
		X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"01",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"97",X"22",X"22",X"22",X"97",X"22",X"22",X"22",X"77",X"22",X"22",X"22",X"79",X"22",
		X"22",X"22",X"7F",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",
		X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",
		X"22",X"22",X"FF",X"22",X"22",X"92",X"FF",X"22",X"2A",X"A9",X"99",X"22",X"AA",X"AA",X"FF",X"22",
		X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"29",X"92",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",
		X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"29",X"92",X"99",X"22",X"22",X"22",X"99",X"22",
		X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"29",X"92",X"99",X"22",X"22",X"22",X"99",X"22",
		X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"29",X"92",X"99",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"29",X"29",X"29",X"22",
		X"92",X"92",X"92",X"22",X"29",X"59",X"29",X"22",X"92",X"55",X"92",X"22",X"29",X"5E",X"29",X"22",
		X"92",X"E5",X"92",X"22",X"29",X"F5",X"29",X"22",X"92",X"F5",X"92",X"22",X"29",X"F5",X"29",X"22",
		X"92",X"FE",X"92",X"22",X"29",X"F5",X"29",X"22",X"92",X"55",X"92",X"22",X"29",X"5E",X"29",X"22",
		X"92",X"55",X"92",X"22",X"29",X"FF",X"29",X"22",X"92",X"95",X"92",X"22",X"29",X"29",X"29",X"22",
		X"92",X"92",X"92",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",
		X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",
		X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",
		X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"05",X"55",X"55",X"00",X"99",X"FF",X"55",
		X"00",X"FF",X"FF",X"FF",X"00",X"FF",X"EE",X"EE",X"00",X"FF",X"99",X"EE",X"00",X"EE",X"9E",X"EE",
		X"00",X"5E",X"E5",X"55",X"99",X"35",X"F9",X"99",X"FF",X"39",X"F9",X"E9",X"FF",X"39",X"F9",X"94",
		X"FF",X"39",X"F9",X"24",X"FF",X"39",X"F9",X"44",X"FF",X"39",X"F9",X"24",X"FE",X"39",X"F9",X"42",
		X"FF",X"39",X"F9",X"24",X"FF",X"39",X"F9",X"42",X"FF",X"39",X"F9",X"24",X"F5",X"39",X"F9",X"22",
		X"F5",X"39",X"F9",X"92",X"FF",X"39",X"F9",X"F9",X"99",X"95",X"F9",X"99",X"05",X"55",X"5F",X"FF",
		X"00",X"5E",X"35",X"55",X"00",X"FF",X"33",X"55",X"00",X"FF",X"55",X"55",X"00",X"FF",X"FF",X"FF",
		X"00",X"5F",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"99",X"09",X"90",X"00",X"55",X"55",X"E0",X"00",
		X"FF",X"FF",X"E0",X"00",X"FF",X"FF",X"E0",X"00",X"F2",X"22",X"E0",X"00",X"22",X"44",X"E0",X"00",
		X"24",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",
		X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",
		X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",
		X"44",X"44",X"E0",X"00",X"44",X"44",X"E0",X"00",X"24",X"24",X"E0",X"00",X"22",X"22",X"E0",X"00",
		X"22",X"22",X"E0",X"00",X"3F",X"FF",X"E0",X"00",X"3F",X"FF",X"E0",X"00",X"FF",X"FF",X"E0",X"00",
		X"FF",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"E0",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"09",X"99",X"55",X"EE",
		X"99",X"44",X"53",X"9E",X"99",X"99",X"59",X"9E",X"99",X"99",X"03",X"9E",X"99",X"99",X"33",X"EE",
		X"44",X"99",X"33",X"E9",X"99",X"99",X"33",X"E5",X"99",X"99",X"39",X"EE",X"AA",X"AA",X"33",X"95",
		X"AA",X"AA",X"93",X"EE",X"AA",X"AA",X"33",X"EE",X"44",X"AA",X"99",X"EE",X"AA",X"AA",X"93",X"9E",
		X"AA",X"AA",X"99",X"9E",X"99",X"AA",X"F9",X"9E",X"99",X"44",X"F9",X"EE",X"09",X"AA",X"FF",X"5E",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",X"00",X"99",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"01",X"00",X"00",X"00",X"99",X"A0",X"00",X"00",X"90",X"A0",X"00",X"06",X"90",X"A0",X"00",
		X"44",X"99",X"AC",X"00",X"46",X"09",X"00",X"00",X"46",X"90",X"00",X"00",X"44",X"99",X"0F",X"00",
		X"06",X"01",X"00",X"00",X"00",X"CA",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"0A",X"00",
		X"44",X"99",X"E0",X"00",X"44",X"90",X"00",X"00",X"44",X"09",X"90",X"00",X"44",X"99",X"A0",X"00",
		X"00",X"90",X"A0",X"00",X"00",X"90",X"A0",X"00",X"00",X"99",X"A0",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"0E",X"00",X"00",X"FE",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0B",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9A",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"50",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"F0",X"A0",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"50",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"9A",X"00",X"00",X"50",X"A0",X"00",
		X"00",X"00",X"A5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"C9",X"99",X"99",X"00",
		X"BC",X"9C",X"99",X"00",X"B6",X"C0",X"CC",X"91",X"AA",X"BE",X"BE",X"10",X"AC",X"9B",X"90",X"91",
		X"AA",X"9B",X"EC",X"11",X"BE",X"9B",X"BE",X"11",X"EB",X"95",X"EB",X"11",X"BE",X"9B",X"BB",X"51",
		X"BB",X"95",X"BB",X"19",X"EE",X"9B",X"BB",X"51",X"5F",X"9F",X"BB",X"59",X"BB",X"9B",X"BB",X"51",
		X"BB",X"9F",X"BB",X"19",X"BB",X"9F",X"BB",X"51",X"6F",X"9F",X"FB",X"11",X"B6",X"9F",X"BF",X"11",
		X"9B",X"9B",X"F9",X"11",X"C9",X"BB",X"BB",X"91",X"BB",X"BB",X"BB",X"10",X"B6",X"C0",X"CC",X"01",
		X"BC",X"9C",X"99",X"00",X"C9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",
		X"99",X"99",X"99",X"00",X"E9",X"99",X"99",X"00",X"E9",X"09",X"59",X"00",X"17",X"99",X"59",X"90",
		X"17",X"99",X"22",X"99",X"19",X"A9",X"D2",X"99",X"99",X"77",X"9E",X"10",X"50",X"D7",X"A9",X"00",
		X"9E",X"7D",X"A9",X"99",X"E9",X"77",X"A9",X"FE",X"E9",X"77",X"A9",X"99",X"5E",X"77",X"AE",X"FE",
		X"59",X"77",X"AE",X"00",X"99",X"77",X"EE",X"10",X"19",X"70",X"D2",X"00",X"17",X"00",X"22",X"00",
		X"16",X"00",X"50",X"00",X"E9",X"00",X"50",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"3E",X"99",X"00",
		X"99",X"EE",X"99",X"00",X"99",X"99",X"99",X"00",X"FF",X"FF",X"99",X"00",X"99",X"99",X"AA",X"00",
		X"A7",X"A7",X"AA",X"00",X"AA",X"AA",X"A9",X"00",X"AA",X"AA",X"95",X"00",X"AA",X"AA",X"99",X"00",
		X"A9",X"AA",X"99",X"00",X"A4",X"AA",X"99",X"00",X"AA",X"AA",X"99",X"00",X"AA",X"AA",X"99",X"00",
		X"AA",X"AA",X"99",X"00",X"AA",X"AA",X"99",X"00",X"A9",X"AA",X"99",X"00",X"A4",X"AA",X"99",X"00",
		X"EA",X"AA",X"99",X"00",X"AE",X"AA",X"05",X"00",X"EE",X"AE",X"A0",X"00",X"EE",X"E5",X"AA",X"00",
		X"99",X"99",X"AA",X"00",X"FF",X"FF",X"99",X"00",X"99",X"99",X"99",X"00",X"D9",X"EE",X"99",X"00",
		X"00",X"3E",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",
		X"E3",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"EA",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"39",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"10",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"61",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"09",X"09",X"90",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"9A",X"AE",X"99",X"5E",X"6E",X"AA",X"99",X"EE",X"6E",X"A9",X"AE",X"99",
		X"6A",X"9A",X"9A",X"9A",X"3A",X"A9",X"FF",X"F9",X"99",X"99",X"9A",X"9A",X"99",X"99",X"99",X"99",
		X"FF",X"9F",X"7A",X"7A",X"F9",X"9F",X"AE",X"AE",X"99",X"FF",X"EA",X"EA",X"99",X"F9",X"AE",X"AE",
		X"FF",X"F9",X"EA",X"EA",X"99",X"99",X"EE",X"AE",X"99",X"99",X"EE",X"EA",X"FF",X"99",X"5E",X"AE",
		X"99",X"F9",X"EE",X"EA",X"99",X"F9",X"5E",X"AE",X"F9",X"FF",X"E5",X"EA",X"FF",X"9F",X"65",X"55",
		X"99",X"9F",X"AA",X"AA",X"99",X"99",X"DD",X"DD",X"39",X"A9",X"FF",X"FD",X"6E",X"AB",X"DD",X"DD",
		X"6E",X"EA",X"AA",X"AA",X"6E",X"AE",X"EE",X"E5",X"0A",X"EE",X"09",X"EE",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"FF",X"91",X"11",X"11",X"5F",X"92",X"11",X"11",X"BF",X"92",X"11",X"11",X"BF",X"92",
		X"11",X"11",X"BF",X"99",X"11",X"99",X"BF",X"99",X"12",X"22",X"BF",X"F9",X"22",X"21",X"AA",X"F9",
		X"19",X"11",X"99",X"F9",X"11",X"21",X"99",X"F9",X"11",X"21",X"FF",X"F9",X"11",X"29",X"BB",X"F9",
		X"11",X"91",X"BB",X"F9",X"11",X"11",X"BB",X"FF",X"11",X"11",X"BB",X"5F",X"12",X"22",X"BB",X"5F",
		X"11",X"11",X"AA",X"5F",X"11",X"91",X"99",X"5F",X"11",X"11",X"99",X"5F",X"91",X"11",X"FF",X"FF",
		X"91",X"11",X"55",X"55",X"91",X"11",X"19",X"99",X"00",X"22",X"22",X"22",X"09",X"11",X"11",X"21",
		X"09",X"11",X"11",X"11",X"09",X"11",X"11",X"22",X"09",X"11",X"11",X"22",X"00",X"19",X"11",X"99",
		X"09",X"91",X"99",X"99",X"09",X"00",X"00",X"00",X"09",X"00",X"EE",X"EE",X"09",X"99",X"99",X"99",
		X"99",X"22",X"29",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"29",X"29",X"22",X"22",X"92",X"99",X"99",
		X"29",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"33",X"33",X"33",X"33",X"93",X"33",X"99",X"92",
		X"33",X"33",X"33",X"33",X"33",X"11",X"33",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"11",X"11",X"22",X"11",X"22",X"22",X"22",X"22",
		X"19",X"11",X"91",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"91",X"91",X"91",X"11",X"19",X"92",X"11",X"22",X"19",X"99",X"91",X"11",X"22",X"99",X"92",
		X"09",X"99",X"99",X"99",X"09",X"33",X"EE",X"EE",X"09",X"33",X"33",X"33",X"09",X"91",X"99",X"99",
		X"00",X"19",X"22",X"22",X"09",X"22",X"22",X"22",X"09",X"22",X"22",X"22",X"09",X"22",X"99",X"22",
		X"09",X"22",X"99",X"22",X"00",X"22",X"99",X"99",X"92",X"22",X"99",X"11",X"92",X"22",X"99",X"22",
		X"92",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"39",X"22",X"29",X"22",X"EE",X"99",
		X"11",X"22",X"EE",X"22",X"22",X"22",X"E2",X"22",X"22",X"22",X"52",X"22",X"22",X"22",X"22",X"22",
		X"29",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"92",X"29",X"92",X"22",X"29",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"F5",X"90",X"00",X"11",X"F5",X"00",X"00",X"11",X"F5",X"00",X"00",X"11",X"F5",X"00",X"00",
		X"11",X"35",X"90",X"00",X"11",X"35",X"00",X"00",X"11",X"F5",X"00",X"00",X"22",X"35",X"00",X"00",
		X"22",X"95",X"90",X"00",X"99",X"95",X"00",X"00",X"11",X"95",X"00",X"00",X"11",X"95",X"00",X"00",
		X"11",X"95",X"90",X"00",X"11",X"95",X"00",X"00",X"11",X"9F",X"00",X"00",X"21",X"9F",X"55",X"00",
		X"19",X"29",X"55",X"00",X"11",X"19",X"5F",X"00",X"11",X"19",X"5F",X"00",X"22",X"19",X"5F",X"00",
		X"22",X"12",X"5F",X"00",X"22",X"12",X"5F",X"00",X"22",X"19",X"5F",X"00",X"22",X"29",X"5F",X"00",
		X"99",X"11",X"5F",X"00",X"11",X"11",X"50",X"00",X"11",X"11",X"00",X"00",X"19",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"99",X"99",X"00",X"00",
		X"29",X"35",X"00",X"00",X"22",X"35",X"00",X"00",X"22",X"35",X"00",X"00",X"22",X"35",X"90",X"00",
		X"22",X"35",X"00",X"00",X"22",X"35",X"00",X"00",X"92",X"35",X"00",X"00",X"22",X"35",X"90",X"00",
		X"29",X"35",X"00",X"00",X"22",X"F5",X"00",X"00",X"22",X"F5",X"00",X"00",X"22",X"F5",X"90",X"00",
		X"22",X"F5",X"00",X"00",X"22",X"35",X"00",X"00",X"33",X"35",X"00",X"00",X"39",X"35",X"90",X"00",
		X"33",X"35",X"00",X"00",X"33",X"35",X"00",X"00",X"11",X"35",X"00",X"00",X"11",X"35",X"90",X"00",
		X"11",X"35",X"00",X"00",X"11",X"F5",X"00",X"00",X"21",X"F5",X"00",X"00",X"11",X"F5",X"90",X"00",
		X"11",X"F5",X"00",X"00",X"11",X"35",X"00",X"00",X"11",X"35",X"00",X"00",X"11",X"35",X"90",X"00",
		X"11",X"35",X"00",X"00",X"11",X"35",X"00",X"00",X"11",X"35",X"00",X"00",X"22",X"35",X"90",X"00",
		X"99",X"99",X"00",X"00",X"E3",X"EE",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"99",X"00",X"00",
		X"12",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"50",X"00",X"22",X"2F",X"5F",X"00",
		X"22",X"29",X"5F",X"00",X"99",X"29",X"5F",X"00",X"11",X"22",X"5F",X"00",X"22",X"22",X"5F",X"00",
		X"22",X"29",X"53",X"00",X"22",X"29",X"3F",X"00",X"99",X"29",X"5F",X"00",X"22",X"F9",X"55",X"00",
		X"22",X"9F",X"55",X"00",X"22",X"9F",X"00",X"00",X"22",X"95",X"00",X"00",X"22",X"95",X"90",X"00",
		X"22",X"25",X"00",X"00",X"22",X"95",X"00",X"00",X"22",X"95",X"00",X"00",X"22",X"F5",X"90",X"00",
		X"33",X"F5",X"00",X"00",X"33",X"F5",X"00",X"00",X"33",X"F5",X"00",X"00",X"92",X"F5",X"90",X"00",
		X"22",X"F5",X"00",X"00",X"22",X"F5",X"00",X"00",X"22",X"F5",X"00",X"00",X"22",X"F5",X"90",X"00",
		X"00",X"09",X"00",X"00",X"00",X"90",X"99",X"90",X"00",X"99",X"11",X"09",X"09",X"55",X"11",X"90",
		X"00",X"55",X"19",X"09",X"99",X"55",X"19",X"99",X"55",X"55",X"19",X"55",X"55",X"55",X"99",X"55",
		X"55",X"33",X"99",X"33",X"55",X"47",X"77",X"33",X"11",X"93",X"39",X"39",X"44",X"33",X"BB",X"41",
		X"55",X"33",X"99",X"95",X"11",X"55",X"99",X"55",X"15",X"55",X"33",X"55",X"55",X"5A",X"11",X"55",
		X"FF",X"5A",X"77",X"55",X"1F",X"55",X"55",X"55",X"11",X"55",X"99",X"F5",X"55",X"55",X"99",X"95",
		X"44",X"FF",X"BB",X"11",X"11",X"11",X"FF",X"FF",X"55",X"41",X"11",X"F5",X"55",X"55",X"99",X"55",
		X"F5",X"55",X"99",X"5F",X"F5",X"55",X"19",X"F0",X"00",X"55",X"19",X"00",X"00",X"FF",X"19",X"00",
		X"00",X"FF",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",X"E9",X"FF",X"00",X"00",
		X"33",X"99",X"00",X"00",X"55",X"39",X"00",X"00",X"59",X"95",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"90",X"00",X"00",
		X"F9",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"FF",X"5F",X"00",X"00",X"FF",X"09",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"60",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"09",X"00",X"00",X"99",X"66",X"60",X"00",X"FF",X"99",X"16",X"00",X"E9",X"FF",X"00",X"00",
		X"33",X"99",X"00",X"00",X"55",X"39",X"00",X"00",X"59",X"95",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"90",X"00",X"00",
		X"F9",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"FF",X"5F",X"00",X"00",X"FF",X"09",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"90",X"06",X"00",X"99",X"F6",X"00",X"00",X"FF",X"01",X"00",X"00",
		X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",X"E9",X"FF",X"00",X"00",
		X"33",X"99",X"00",X"00",X"55",X"39",X"00",X"00",X"59",X"95",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"90",X"00",X"00",
		X"F9",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"FF",X"5F",X"00",X"00",X"FF",X"09",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"F0",X"60",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"61",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"09",X"00",X"00",X"99",X"99",X"00",X"09",X"22",X"22",X"00",X"92",X"11",X"11",
		X"00",X"21",X"77",X"11",X"00",X"11",X"22",X"22",X"00",X"77",X"29",X"29",X"00",X"22",X"92",X"92",
		X"00",X"29",X"99",X"29",X"01",X"22",X"44",X"99",X"11",X"44",X"94",X"49",X"1C",X"44",X"49",X"29",
		X"CC",X"44",X"99",X"29",X"C9",X"44",X"22",X"29",X"92",X"44",X"22",X"29",X"92",X"41",X"62",X"29",
		X"99",X"16",X"96",X"29",X"92",X"1F",X"26",X"29",X"99",X"76",X"96",X"99",X"92",X"7F",X"62",X"99",
		X"99",X"47",X"24",X"99",X"C9",X"44",X"44",X"29",X"12",X"44",X"44",X"29",X"C1",X"44",X"44",X"49",
		X"1C",X"46",X"44",X"22",X"11",X"99",X"92",X"22",X"07",X"92",X"29",X"29",X"00",X"99",X"92",X"99",
		X"00",X"22",X"99",X"21",X"00",X"11",X"22",X"11",X"00",X"11",X"11",X"11",X"00",X"06",X"72",X"20",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"22",X"99",X"00",X"00",
		X"11",X"22",X"90",X"00",X"11",X"11",X"09",X"00",X"22",X"21",X"90",X"00",X"92",X"22",X"29",X"00",
		X"99",X"29",X"22",X"00",X"77",X"92",X"12",X"00",X"77",X"99",X"12",X"00",X"27",X"22",X"11",X"00",
		X"77",X"29",X"11",X"00",X"22",X"F2",X"21",X"00",X"77",X"29",X"11",X"00",X"22",X"F2",X"21",X"00",
		X"22",X"29",X"10",X"00",X"22",X"F2",X"21",X"00",X"22",X"29",X"11",X"00",X"22",X"F2",X"21",X"00",
		X"22",X"29",X"11",X"00",X"99",X"F2",X"11",X"00",X"92",X"99",X"12",X"00",X"49",X"22",X"10",X"00",
		X"22",X"92",X"00",X"00",X"22",X"29",X"00",X"00",X"92",X"92",X"00",X"00",X"99",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"12",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"50",X"55",X"00",X"00",X"55",X"55",X"00",X"00",
		X"5F",X"5F",X"00",X"00",X"05",X"5F",X"00",X"00",X"50",X"05",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"05",X"00",X"05",X"55",X"5F",X"50",
		X"5F",X"05",X"5F",X"00",X"05",X"50",X"05",X"00",X"50",X"05",X"55",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"50",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",
		X"0F",X"55",X"00",X"00",X"05",X"55",X"00",X"00",X"50",X"55",X"00",X"00",X"05",X"05",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"50",X"00",X"00",
		X"F1",X"55",X"00",X"00",X"1F",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"51",X"55",X"00",X"00",
		X"55",X"55",X"00",X"00",X"F5",X"55",X"00",X"00",X"FF",X"15",X"50",X"00",X"FF",X"11",X"55",X"00",
		X"FF",X"11",X"55",X"00",X"FF",X"11",X"55",X"00",X"1F",X"31",X"55",X"00",X"1F",X"53",X"55",X"00",
		X"1F",X"55",X"11",X"00",X"1F",X"99",X"11",X"00",X"11",X"99",X"11",X"00",X"11",X"BB",X"19",X"90",
		X"11",X"99",X"99",X"00",X"11",X"99",X"95",X"00",X"51",X"99",X"12",X"09",X"51",X"99",X"12",X"00",
		X"55",X"99",X"11",X"09",X"55",X"91",X"F1",X"00",X"55",X"B9",X"B1",X"00",X"55",X"BB",X"91",X"00",
		X"55",X"FB",X"99",X"09",X"55",X"FB",X"99",X"00",X"F5",X"1F",X"95",X"09",X"05",X"11",X"5F",X"90",
		X"55",X"35",X"99",X"00",X"95",X"35",X"99",X"90",X"0F",X"33",X"19",X"96",X"00",X"13",X"11",X"96",
		X"00",X"11",X"31",X"00",X"90",X"51",X"31",X"90",X"09",X"F1",X"F3",X"99",X"90",X"FF",X"99",X"99",
		X"00",X"FF",X"FF",X"F6",X"00",X"F9",X"99",X"00",X"00",X"F9",X"9F",X"06",X"00",X"F9",X"FF",X"00",
		X"00",X"F9",X"9F",X"F0",X"00",X"F9",X"3F",X"00",X"00",X"F9",X"3F",X"90",X"00",X"0F",X"13",X"00",
		X"00",X"0F",X"11",X"09",X"00",X"0F",X"F1",X"00",X"00",X"00",X"F2",X"90",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"90",X"00",X"99",X"59",X"D9",X"00",X"00",X"9B",X"B9",X"00",X"00",X"99",X"90",
		X"00",X"99",X"00",X"00",X"00",X"BA",X"00",X"00",X"09",X"AB",X"90",X"00",X"94",X"BA",X"99",X"00",
		X"99",X"9B",X"D9",X"00",X"D9",X"44",X"99",X"00",X"D9",X"F4",X"BA",X"BB",X"99",X"F4",X"BB",X"BB",
		X"9B",X"F4",X"BB",X"99",X"BB",X"F4",X"BB",X"B5",X"BB",X"F4",X"BB",X"99",X"BB",X"94",X"BB",X"FF",
		X"FB",X"F4",X"BB",X"99",X"BF",X"94",X"BB",X"55",X"FB",X"F4",X"BF",X"99",X"AA",X"94",X"FB",X"B5",
		X"BA",X"94",X"BA",X"BB",X"BA",X"44",X"99",X"00",X"BA",X"9B",X"AA",X"00",X"A4",X"BB",X"A9",X"00",
		X"0A",X"BA",X"90",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"99",X"90",
		X"00",X"00",X"9D",X"D9",X"00",X"99",X"59",X"B9",X"00",X"00",X"99",X"B9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",X"AE",X"00",X"00",
		X"DB",X"DA",X"00",X"00",X"BD",X"BD",X"DA",X"00",X"BB",X"BB",X"BB",X"90",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"5B",X"A0",X"BB",X"BB",X"BA",X"00",X"DB",X"BA",X"00",X"00",X"AA",X"AE",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"00",X"00",X"02",X"F4",X"00",X"00",X"22",X"F4",X"00",X"00",X"22",X"FF",X"00",X"00",
		X"22",X"FF",X"00",X"00",X"22",X"9F",X"00",X"00",X"22",X"99",X"90",X"00",X"99",X"44",X"D9",X"00",
		X"BA",X"FF",X"D9",X"90",X"BB",X"FF",X"DD",X"99",X"BB",X"FF",X"DD",X"D9",X"BB",X"FF",X"9D",X"DD",
		X"BB",X"F9",X"B9",X"9D",X"AB",X"9F",X"BB",X"9B",X"9B",X"99",X"BB",X"90",X"0B",X"94",X"BB",X"00",
		X"09",X"94",X"BB",X"90",X"00",X"4F",X"BB",X"90",X"00",X"B9",X"BB",X"B9",X"99",X"AA",X"BB",X"BB",
		X"00",X"AA",X"B9",X"BB",X"99",X"AA",X"B9",X"B9",X"09",X"AA",X"99",X"99",X"00",X"00",X"99",X"9F",
		X"00",X"00",X"99",X"9F",X"00",X"00",X"99",X"5F",X"00",X"00",X"99",X"55",X"00",X"90",X"99",X"D5",
		X"00",X"0F",X"99",X"DD",X"00",X"0B",X"90",X"0D",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"DE",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"D0",X"00",X"00",
		X"BB",X"BD",X"0D",X"00",X"DD",X"BB",X"0D",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"BF",X"0A",X"00",X"00",X"BB",X"0A",X"00",X"00",X"DB",X"AA",X"00",X"00",X"00",X"DA",X"00",
		X"00",X"00",X"BD",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"DF",X"00",
		X"00",X"00",X"BD",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"D9",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"BB",X"90",X"00",X"00",X"BB",X"99",X"00",X"00",X"BA",X"99",X"00",X"00",
		X"B4",X"99",X"00",X"00",X"44",X"9D",X"00",X"00",X"4F",X"99",X"00",X"00",X"9F",X"9D",X"90",X"00",
		X"9F",X"99",X"90",X"00",X"99",X"9D",X"99",X"00",X"9F",X"99",X"99",X"00",X"99",X"9D",X"09",X"00",
		X"9F",X"B9",X"00",X"00",X"99",X"B9",X"00",X"00",X"44",X"BB",X"0D",X"00",X"44",X"BB",X"0B",X"00",
		X"4F",X"BB",X"0B",X"00",X"9F",X"BB",X"0B",X"00",X"99",X"BA",X"99",X"00",X"A9",X"BB",X"99",X"00",
		X"A9",X"BA",X"99",X"00",X"A9",X"BB",X"99",X"00",X"99",X"B9",X"99",X"00",X"99",X"99",X"00",X"00",
		X"99",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"B9",X"00",X"00",
		X"00",X"B9",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"90",X"0A",X"00",X"00",
		X"99",X"00",X"A0",X"00",X"D9",X"00",X"A0",X"00",X"DD",X"00",X"D0",X"00",X"BD",X"00",X"DD",X"00",
		X"BD",X"00",X"BA",X"00",X"0B",X"00",X"BD",X"00",X"0B",X"00",X"BD",X"00",X"00",X"00",X"FB",X"DD",
		X"00",X"00",X"55",X"DD",X"00",X"00",X"BF",X"DD",X"00",X"00",X"DB",X"0D",X"00",X"00",X"DB",X"0B",
		X"00",X"00",X"0D",X"BB",X"00",X"00",X"0D",X"A9",X"00",X"00",X"0D",X"A9",X"00",X"00",X"00",X"A9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",X"A0",X"00",X"00",X"A9",X"A0",X"00",X"00",X"AA",X"A0",
		X"00",X"B5",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"DB",X"00",X"00",X"00",X"B5",X"00",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"D5",X"00",X"00",
		X"00",X"DB",X"00",X"00",X"00",X"D5",X"00",X"00",X"00",X"DB",X"00",X"00",X"00",X"D5",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"0A",X"BD",X"A0",X"00",X"0A",X"BD",X"AB",X"00",X"0A",X"BD",X"AB",X"00",
		X"0A",X"BA",X"BB",X"00",X"0A",X"0A",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"90",X"00",
		X"00",X"99",X"D9",X"00",X"00",X"AF",X"DD",X"00",X"00",X"AF",X"D9",X"00",X"00",X"FB",X"99",X"00",
		X"99",X"44",X"44",X"00",X"00",X"49",X"FB",X"00",X"00",X"49",X"BF",X"00",X"00",X"99",X"F4",X"00",
		X"00",X"9F",X"49",X"00",X"00",X"99",X"9D",X"00",X"00",X"99",X"D9",X"00",X"00",X"44",X"9D",X"00",
		X"00",X"FB",X"DD",X"00",X"99",X"BF",X"DD",X"00",X"00",X"FB",X"DD",X"00",X"00",X"BB",X"DD",X"00",
		X"00",X"FB",X"DD",X"00",X"00",X"BB",X"D9",X"00",X"00",X"BB",X"99",X"00",X"00",X"BB",X"90",X"00",
		X"00",X"BB",X"90",X"00",X"00",X"BB",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"B5",X"99",X"00",X"99",X"59",X"99",X"00",X"99",X"59",X"99",X"00",X"99",X"59",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"00",X"06",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"64",X"00",
		X"00",X"40",X"66",X"00",X"00",X"64",X"66",X"00",X"04",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"46",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"04",X"60",X"00",
		X"04",X"46",X"40",X"00",X"46",X"66",X"00",X"00",X"00",X"66",X"40",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"40",X"00",X"04",X"66",X"60",X"00",
		X"00",X"64",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"06",X"40",X"00",X"00",X"06",X"60",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"06",X"00",
		X"00",X"40",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"06",X"00",X"00",
		X"00",X"06",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"40",X"00",X"66",X"00",X"66",X"00",
		X"06",X"40",X"66",X"00",X"00",X"64",X"64",X"00",X"04",X"06",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"40",X"66",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"60",X"00",X"60",X"04",X"60",X"00",
		X"64",X"46",X"40",X"00",X"40",X"66",X"00",X"00",X"00",X"66",X"40",X"00",X"00",X"40",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"40",X"00",X"04",X"66",X"66",X"00",
		X"06",X"64",X"66",X"00",X"66",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"06",X"40",X"00",X"00",X"06",X"60",X"00",X"00",X"60",X"60",X"00",X"00",X"00",X"06",X"00",
		X"00",X"40",X"00",X"00",X"00",X"66",X"04",X"00",X"04",X"66",X"40",X"00",X"06",X"66",X"00",X"00",
		X"00",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"40",X"00",X"66",X"04",X"66",X"00",
		X"06",X"40",X"66",X"00",X"00",X"66",X"64",X"00",X"04",X"66",X"46",X"00",X"00",X"60",X"66",X"00",
		X"00",X"40",X"66",X"00",X"06",X"00",X"00",X"00",X"40",X"66",X"60",X"00",X"60",X"64",X"60",X"00",
		X"04",X"46",X"40",X"00",X"40",X"66",X"00",X"00",X"66",X"66",X"40",X"00",X"00",X"46",X"60",X"00",
		X"00",X"66",X"66",X"00",X"04",X"66",X"60",X"00",X"66",X"66",X"40",X"00",X"66",X"66",X"66",X"00",
		X"66",X"64",X"64",X"00",X"66",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"00",X"06",X"66",X"00",
		X"00",X"00",X"40",X"00",X"06",X"60",X"60",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"40",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"40",X"00",X"66",X"04",X"66",X"00",
		X"64",X"40",X"66",X"00",X"00",X"06",X"64",X"00",X"04",X"66",X"46",X"44",X"00",X"60",X"66",X"60",
		X"60",X"40",X"66",X"00",X"06",X"00",X"66",X"00",X"46",X"00",X"60",X"00",X"00",X"00",X"60",X"00",
		X"46",X"06",X"40",X"00",X"66",X"66",X"00",X"00",X"66",X"00",X"40",X"00",X"00",X"40",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"06",X"60",X"00",X"00",X"66",X"40",X"00",X"66",X"60",X"66",X"00",
		X"66",X"04",X"64",X"00",X"66",X"00",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"40",X"66",X"00",
		X"60",X"00",X"66",X"00",X"06",X"E0",X"60",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"0A",X"A0",X"00",
		X"0A",X"A0",X"00",X"00",X"00",X"0A",X"0F",X"00",X"A0",X"A0",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"A0",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"0A",X"00",X"A0",X"00",
		X"A0",X"0A",X"00",X"00",X"FF",X"A0",X"A0",X"00",X"00",X"0A",X"0A",X"00",X"0F",X"0F",X"A0",X"00",
		X"00",X"F0",X"0A",X"00",X"F0",X"0F",X"F0",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"0A",X"0A",X"00",X"A0",X"A0",X"A0",X"0A",X"00",
		X"00",X"0A",X"00",X"00",X"AA",X"00",X"F0",X"00",X"0F",X"0F",X"0F",X"00",X"F0",X"A0",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"A0",X"0A",X"00",X"00",X"00",X"00",X"0A",X"00",X"0F",X"A0",X"A0",X"00",
		X"00",X"FA",X"00",X"00",X"0F",X"00",X"A0",X"00",X"00",X"0F",X"0A",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"FF",X"FF",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"FF",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"FF",X"F0",X"00",
		X"00",X"F0",X"0F",X"00",X"00",X"FF",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"0F",X"FF",X"FF",X"00",
		X"F0",X"FF",X"00",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"0F",X"0F",X"F0",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"F0",X"F0",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"F0",X"0F",X"00",X"00",X"0F",X"00",X"00",X"F0",X"F0",X"F0",X"00",X"0F",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"39",X"00",X"00",X"93",X"B3",X"00",X"00",X"BB",X"5B",X"39",X"00",
		X"BB",X"5F",X"93",X"00",X"93",X"B3",X"00",X"00",X"09",X"39",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"39",X"00",X"00",X"93",X"B3",X"00",X"00",X"B5",X"55",X"39",X"00",
		X"BB",X"5F",X"93",X"00",X"93",X"B3",X"00",X"00",X"09",X"39",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"93",X"00",X"00",X"30",X"30",X"00",X"00",X"05",X"03",X"50",X"00",
		X"05",X"00",X"0F",X"50",X"30",X"30",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"93",X"00",X"00",X"30",X"30",X"00",X"00",X"05",X"03",X"05",X"00",
		X"05",X"00",X"00",X"05",X"30",X"30",X"F0",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"00",X"9D",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"DD",X"99",X"99",X"00",X"9D",X"99",X"99",X"09",X"D9",X"99",X"EE",X"99",X"EE",X"99",X"99",
		X"DD",X"59",X"E5",X"55",X"99",X"39",X"B9",X"99",X"DD",X"99",X"59",X"E9",X"99",X"99",X"B9",X"9A",
		X"DD",X"99",X"59",X"AB",X"99",X"99",X"B9",X"BA",X"DD",X"99",X"59",X"AB",X"99",X"EE",X"B9",X"BA",
		X"AA",X"BB",X"B9",X"AB",X"AB",X"99",X"B9",X"BA",X"BA",X"99",X"59",X"AB",X"AB",X"99",X"B5",X"9A",
		X"BA",X"99",X"59",X"9A",X"AB",X"99",X"B9",X"F9",X"BA",X"99",X"59",X"99",X"AB",X"B9",X"55",X"55",
		X"BA",X"5B",X"95",X"55",X"0B",X"A5",X"99",X"55",X"00",X"BA",X"BA",X"AA",X"00",X"AB",X"AB",X"BB",
		X"00",X"BA",X"BA",X"AA",X"00",X"AB",X"AB",X"BB",X"00",X"BA",X"BA",X"0A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"99",X"D9",X"90",X"00",X"9D",X"9D",X"90",X"00",
		X"DD",X"DB",X"90",X"00",X"9D",X"99",X"90",X"00",X"EB",X"55",X"90",X"00",X"ED",X"DD",X"90",X"00",
		X"EB",X"BB",X"90",X"00",X"ED",X"DD",X"90",X"00",X"EB",X"BB",X"90",X"00",X"ED",X"DD",X"90",X"00",
		X"EB",X"BB",X"90",X"00",X"EB",X"DB",X"90",X"00",X"EB",X"BB",X"90",X"00",X"EB",X"BB",X"90",X"00",
		X"EB",X"BA",X"90",X"00",X"EB",X"BB",X"90",X"00",X"EB",X"AB",X"90",X"00",X"EB",X"BB",X"90",X"00",
		X"EA",X"AA",X"90",X"00",X"EB",X"BB",X"90",X"00",X"EA",X"AA",X"90",X"00",X"EB",X"BB",X"90",X"00",
		X"EA",X"55",X"90",X"00",X"5B",X"B9",X"90",X"00",X"AA",X"AA",X"90",X"00",X"BA",X"AA",X"90",X"00",
		X"AA",X"AA",X"A0",X"00",X"AB",X"AA",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"9A",X"90",X"00",X"9B",X"AB",X"90",X"00",X"9D",X"BD",X"90",X"00",X"9B",X"BB",X"90",
		X"00",X"5B",X"5B",X"90",X"00",X"9A",X"BA",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"9A",X"BA",X"90",
		X"00",X"AB",X"AB",X"90",X"00",X"9B",X"BB",X"90",X"00",X"B5",X"B5",X"90",X"00",X"9B",X"AB",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"F0",X"F0",X"0F",X"00",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"0F",X"00",X"0F",X"5F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"00",X"F0",X"FF",X"F0",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"0F",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"0F",X"F0",X"0F",X"00",X"FF",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",
		X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"50",X"0F",X"0F",
		X"00",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AF",X"00",X"00",X"99",X"5A",X"00",X"00",X"99",X"95",X"00",X"00",X"95",X"55",X"00",
		X"00",X"95",X"51",X"99",X"99",X"55",X"51",X"55",X"09",X"55",X"11",X"33",X"99",X"55",X"11",X"33",
		X"00",X"33",X"77",X"77",X"09",X"44",X"39",X"93",X"09",X"39",X"BB",X"33",X"99",X"33",X"B9",X"D9",
		X"9F",X"53",X"99",X"D9",X"89",X"33",X"99",X"D9",X"01",X"35",X"99",X"D9",X"09",X"35",X"99",X"D9",
		X"99",X"33",X"99",X"D9",X"89",X"F3",X"91",X"D9",X"59",X"FF",X"91",X"39",X"99",X"99",X"95",X"33",
		X"99",X"11",X"9F",X"F5",X"99",X"55",X"99",X"11",X"09",X"55",X"11",X"55",X"00",X"95",X"11",X"55",
		X"00",X"99",X"51",X"FF",X"00",X"99",X"51",X"00",X"00",X"9F",X"55",X"00",X"00",X"98",X"FF",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"09",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"9F",X"00",X"00",X"9F",X"F3",X"00",X"00",
		X"FF",X"33",X"3F",X"00",X"95",X"33",X"00",X"00",X"13",X"03",X"00",X"00",X"93",X"03",X"00",X"00",
		X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",
		X"9F",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"99",X"99",X"00",X"00",X"11",X"11",X"00",X"00",
		X"55",X"FF",X"00",X"00",X"99",X"F0",X"0F",X"00",X"99",X"90",X"00",X"00",X"F9",X"99",X"0F",X"00",
		X"0F",X"99",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"FF",X"00",X"0F",X"0F",X"00",X"00",X"90",X"00",X"00",X"00",X"95",X"50",X"FF",
		X"00",X"99",X"95",X"00",X"09",X"55",X"55",X"55",X"00",X"99",X"51",X"33",X"99",X"95",X"11",X"33",
		X"00",X"33",X"77",X"77",X"00",X"44",X"33",X"99",X"00",X"73",X"AB",X"33",X"85",X"33",X"BB",X"9D",
		X"08",X"55",X"B9",X"9D",X"88",X"53",X"99",X"DD",X"00",X"33",X"99",X"DD",X"00",X"53",X"99",X"DD",
		X"09",X"F3",X"99",X"DD",X"08",X"FF",X"B9",X"9D",X"05",X"FF",X"99",X"93",X"09",X"1F",X"99",X"39",
		X"89",X"11",X"99",X"99",X"99",X"55",X"99",X"99",X"00",X"55",X"99",X"55",X"00",X"95",X"99",X"55",
		X"00",X"99",X"99",X"0F",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",X"00",X"09",X"9F",X"00",
		X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"30",X"00",
		X"FF",X"00",X"03",X"00",X"59",X"00",X"30",X"00",X"11",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"F3",X"00",X"F0",X"00",X"F3",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"F0",X"F0",X"00",
		X"F9",X"00",X"F0",X"00",X"FF",X"0F",X"00",X"00",X"99",X"0F",X"F0",X"00",X"11",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"99",X"00",X"00",
		X"F0",X"F9",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"0F",X"0F",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"FF",X"0F",X"0F",X"0F",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"0F",X"55",X"51",X"30",
		X"00",X"55",X"11",X"33",X"00",X"33",X"77",X"77",X"00",X"44",X"33",X"99",X"00",X"73",X"AB",X"03",
		X"89",X"33",X"BB",X"0D",X"09",X"55",X"B9",X"0D",X"88",X"53",X"99",X"0D",X"00",X"33",X"99",X"DD",
		X"00",X"53",X"99",X"DD",X"09",X"F3",X"99",X"DD",X"08",X"FF",X"B9",X"9D",X"05",X"FF",X"99",X"93",
		X"09",X"1F",X"99",X"39",X"89",X"91",X"FF",X"99",X"99",X"55",X"55",X"99",X"00",X"55",X"55",X"11",
		X"00",X"99",X"55",X"11",X"00",X"99",X"55",X"55",X"00",X"99",X"55",X"55",X"00",X"99",X"59",X"99",
		X"00",X"09",X"9F",X"99",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"F0",X"F0",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"09",X"0F",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"F0",X"F0",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"09",X"55",X"00",X"0F",X"95",X"55",X"50",
		X"0F",X"55",X"31",X"00",X"00",X"53",X"77",X"00",X"0F",X"14",X"33",X"00",X"F0",X"47",X"33",X"00",
		X"00",X"71",X"3A",X"00",X"0F",X"55",X"AB",X"00",X"F0",X"55",X"A0",X"00",X"00",X"55",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"F0",X"FF",X"9B",X"09",X"0F",X"FF",X"9B",X"00",X"F0",X"11",X"99",X"00",
		X"00",X"00",X"99",X"90",X"00",X"10",X"99",X"00",X"0F",X"00",X"15",X"90",X"00",X"00",X"55",X"10",
		X"0F",X"00",X"55",X"00",X"00",X"00",X"55",X"10",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"11",X"0F",X"F0",X"00",X"11",X"00",X"00",X"00",
		X"15",X"00",X"F0",X"00",X"59",X"0F",X"0F",X"00",X"99",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"09",X"99",X"00",X"00",X"99",X"33",X"09",X"00",X"15",X"FF",X"00",X"00",X"11",X"F5",X"00",X"00",
		X"11",X"55",X"90",X"00",X"51",X"55",X"99",X"00",X"55",X"55",X"99",X"90",X"55",X"11",X"99",X"90",
		X"55",X"11",X"19",X"00",X"55",X"99",X"11",X"00",X"F5",X"99",X"11",X"90",X"FF",X"99",X"11",X"09",
		X"FF",X"99",X"19",X"00",X"FF",X"9B",X"19",X"09",X"1F",X"9B",X"99",X"99",X"11",X"B9",X"B9",X"99",
		X"11",X"B9",X"9B",X"39",X"99",X"B9",X"99",X"99",X"99",X"B9",X"99",X"F9",X"99",X"B9",X"99",X"99",
		X"99",X"19",X"9D",X"99",X"F9",X"11",X"9D",X"99",X"F5",X"11",X"DD",X"90",X"F5",X"11",X"DF",X"00",
		X"FF",X"11",X"D9",X"00",X"99",X"11",X"11",X"00",X"09",X"11",X"55",X"99",X"09",X"11",X"55",X"99",
		X"00",X"21",X"FF",X"99",X"00",X"F1",X"FF",X"90",X"00",X"F1",X"0F",X"90",X"00",X"F1",X"00",X"F9",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"09",X"00",X"FF",X"10",X"99",X"00",
		X"99",X"11",X"FF",X"00",X"09",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"09",X"99",X"00",X"99",X"00",X"99",X"00",X"9F",X"00",X"FF",X"00",X"99",X"F3",X"33",X"00",
		X"99",X"F5",X"55",X"00",X"09",X"59",X"59",X"00",X"11",X"11",X"11",X"00",X"99",X"11",X"99",X"00",
		X"00",X"FF",X"FF",X"00",X"99",X"F9",X"FF",X"00",X"99",X"F9",X"FF",X"00",X"9F",X"F9",X"FF",X"00",
		X"FF",X"F9",X"FF",X"00",X"FF",X"FF",X"FF",X"00",X"99",X"99",X"99",X"00",X"99",X"14",X"11",X"00",
		X"99",X"11",X"FF",X"00",X"99",X"9F",X"F5",X"00",X"99",X"9E",X"00",X"00",X"90",X"99",X"99",X"00",
		X"00",X"F9",X"99",X"00",X"0F",X"0F",X"FF",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"29",X"99",X"99",X"99",
		X"92",X"22",X"22",X"22",X"29",X"22",X"22",X"22",X"92",X"92",X"22",X"22",X"99",X"99",X"99",X"99",
		X"29",X"29",X"22",X"22",X"99",X"92",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"22",X"99",X"99",
		X"32",X"C2",X"99",X"99",X"32",X"22",X"92",X"2C",X"99",X"C2",X"22",X"22",X"CC",X"92",X"9C",X"2C",
		X"22",X"C9",X"99",X"9C",X"2C",X"2C",X"2C",X"92",X"CC",X"C2",X"2C",X"22",X"22",X"C2",X"22",X"CC",
		X"99",X"99",X"22",X"C2",X"00",X"22",X"99",X"99",X"C0",X"22",X"22",X"2C",X"CC",X"22",X"22",X"C2",
		X"C2",X"2C",X"22",X"2C",X"C9",X"22",X"92",X"99",X"99",X"99",X"99",X"99",X"2C",X"22",X"2C",X"33",
		X"2C",X"22",X"C9",X"33",X"C2",X"22",X"C9",X"93",X"C2",X"2C",X"C2",X"33",X"22",X"C2",X"2C",X"33",
		X"99",X"99",X"9F",X"00",X"22",X"22",X"29",X"00",X"22",X"22",X"2F",X"F0",X"99",X"99",X"99",X"00",
		X"22",X"22",X"29",X"2F",X"22",X"22",X"29",X"0F",X"22",X"22",X"29",X"F0",X"99",X"99",X"99",X"FF",
		X"22",X"22",X"99",X"0F",X"22",X"22",X"99",X"00",X"22",X"32",X"99",X"F0",X"99",X"99",X"9F",X"FF",
		X"00",X"0F",X"0F",X"0F",X"99",X"00",X"0F",X"F0",X"92",X"00",X"F0",X"00",X"29",X"90",X"00",X"00",
		X"22",X"20",X"00",X"00",X"99",X"90",X"00",X"00",X"22",X"92",X"00",X"00",X"99",X"29",X"00",X"00",
		X"22",X"22",X"F0",X"00",X"29",X"92",X"00",X"00",X"99",X"99",X"00",X"F0",X"29",X"22",X"00",X"F0",
		X"2C",X"92",X"0F",X"00",X"22",X"22",X"00",X"00",X"29",X"92",X"00",X"F0",X"99",X"92",X"F0",X"00",
		X"92",X"20",X"00",X"00",X"22",X"22",X"00",X"0F",X"22",X"20",X"F0",X"00",X"92",X"92",X"F0",X"F0",
		X"C2",X"92",X"92",X"99",X"2C",X"22",X"22",X"22",X"C2",X"22",X"22",X"C2",X"2C",X"22",X"22",X"2C",
		X"22",X"99",X"22",X"99",X"9C",X"99",X"29",X"22",X"C2",X"99",X"99",X"CC",X"CC",X"99",X"90",X"22",
		X"CC",X"99",X"09",X"22",X"C2",X"99",X"92",X"C2",X"C9",X"99",X"99",X"99",X"C2",X"29",X"22",X"92",
		X"C2",X"22",X"22",X"22",X"C2",X"22",X"22",X"22",X"2C",X"29",X"29",X"C9",X"2C",X"22",X"99",X"32",
		X"CC",X"99",X"22",X"22",X"3C",X"29",X"29",X"29",X"C3",X"22",X"22",X"22",X"33",X"22",X"22",X"92",
		X"93",X"2C",X"99",X"99",X"33",X"9C",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"20",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"2F",X"00",X"00",
		X"99",X"92",X"F0",X"00",X"22",X"90",X"0F",X"F0",X"22",X"22",X"00",X"F0",X"22",X"20",X"F0",X"00",
		X"22",X"22",X"00",X"0F",X"93",X"92",X"00",X"0F",X"22",X"29",X"F0",X"00",X"92",X"92",X"0F",X"00",
		X"22",X"92",X"F0",X"00",X"93",X"22",X"00",X"00",X"29",X"93",X"F0",X"00",X"92",X"92",X"F0",X"00",
		X"92",X"22",X"F0",X"00",X"29",X"92",X"0F",X"00",X"33",X"99",X"0F",X"0F",X"29",X"22",X"F0",X"00",
		X"92",X"22",X"FF",X"0F",X"22",X"20",X"00",X"00",X"92",X"90",X"00",X"F0",X"99",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"0F",X"F0",X"FF",X"00",X"0F",X"00",X"09",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"22",X"00",X"00",X"0F",X"22",X"00",X"0F",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"92",X"0F",X"00",X"00",X"92",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"29",X"99",X"99",X"99",
		X"92",X"22",X"22",X"22",X"29",X"22",X"22",X"22",X"92",X"92",X"22",X"22",X"99",X"99",X"99",X"99",
		X"29",X"29",X"22",X"22",X"99",X"92",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"22",X"99",X"99",
		X"32",X"C2",X"99",X"99",X"32",X"22",X"92",X"2C",X"99",X"C2",X"22",X"22",X"CC",X"92",X"9C",X"2C",
		X"22",X"C9",X"99",X"9C",X"2C",X"2C",X"2C",X"92",X"CC",X"C2",X"2C",X"22",X"22",X"C2",X"22",X"CC",
		X"99",X"99",X"22",X"C2",X"00",X"22",X"99",X"99",X"C0",X"22",X"22",X"2C",X"CC",X"22",X"22",X"C2",
		X"C2",X"2C",X"22",X"2C",X"C9",X"22",X"92",X"99",X"99",X"99",X"99",X"99",X"2C",X"22",X"2C",X"33",
		X"2C",X"22",X"C9",X"33",X"C2",X"22",X"C9",X"93",X"C2",X"2C",X"C2",X"33",X"22",X"C2",X"2C",X"33",
		X"99",X"99",X"99",X"00",X"22",X"22",X"29",X"00",X"22",X"22",X"29",X"00",X"99",X"99",X"99",X"00",
		X"22",X"22",X"29",X"20",X"22",X"22",X"29",X"0F",X"22",X"22",X"29",X"2F",X"99",X"99",X"99",X"20",
		X"22",X"22",X"99",X"0F",X"22",X"22",X"99",X"00",X"22",X"32",X"99",X"0F",X"99",X"99",X"90",X"0F",
		X"00",X"00",X"0F",X"0F",X"99",X"00",X"F0",X"F0",X"92",X"00",X"F0",X"00",X"29",X"99",X"0F",X"00",
		X"22",X"22",X"00",X"0F",X"99",X"92",X"00",X"00",X"22",X"92",X"00",X"F0",X"99",X"29",X"0F",X"00",
		X"22",X"22",X"F0",X"F0",X"29",X"92",X"00",X"00",X"99",X"99",X"00",X"00",X"29",X"22",X"F0",X"00",
		X"2C",X"92",X"00",X"00",X"22",X"22",X"00",X"F0",X"29",X"22",X"00",X"F0",X"99",X"22",X"0F",X"F0",
		X"92",X"20",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"20",X"00",X"00",X"92",X"22",X"00",X"00",
		X"C2",X"92",X"92",X"99",X"2C",X"22",X"22",X"22",X"C2",X"22",X"22",X"C2",X"2C",X"22",X"22",X"2C",
		X"22",X"99",X"22",X"99",X"9C",X"99",X"29",X"22",X"C2",X"99",X"99",X"CC",X"CC",X"99",X"90",X"22",
		X"CC",X"99",X"09",X"22",X"C2",X"99",X"92",X"C2",X"C9",X"99",X"99",X"99",X"C2",X"29",X"22",X"92",
		X"C2",X"22",X"22",X"22",X"C2",X"22",X"22",X"22",X"2C",X"29",X"29",X"C9",X"2C",X"22",X"99",X"32",
		X"CC",X"99",X"22",X"22",X"3C",X"29",X"29",X"29",X"C3",X"22",X"22",X"22",X"33",X"22",X"22",X"92",
		X"93",X"2C",X"99",X"99",X"33",X"9C",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"20",X"00",X"00",X"99",X"22",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"02",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"20",X"00",X"00",
		X"99",X"22",X"0F",X"00",X"22",X"92",X"00",X"00",X"22",X"22",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"22",X"00",X"00",X"93",X"92",X"00",X"00",X"22",X"29",X"00",X"00",X"92",X"92",X"00",X"00",
		X"22",X"92",X"0F",X"00",X"93",X"22",X"00",X"00",X"29",X"93",X"00",X"00",X"92",X"92",X"0F",X"0F",
		X"92",X"22",X"00",X"00",X"29",X"92",X"00",X"00",X"33",X"99",X"00",X"00",X"29",X"22",X"0F",X"00",
		X"92",X"22",X"F0",X"00",X"22",X"20",X"F0",X"00",X"92",X"90",X"0F",X"00",X"99",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"F0",X"00",X"00",X"09",X"0F",X"00",X"00",X"92",X"F0",X"00",
		X"00",X"22",X"F0",X"00",X"00",X"22",X"F0",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"FF",X"00",
		X"00",X"99",X"F0",X"00",X"00",X"92",X"00",X"00",X"00",X"92",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"0A",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"AA",X"00",X"00",X"9A",X"A7",X"A0",X"00",
		X"9A",X"AE",X"9A",X"00",X"93",X"EA",X"99",X"AA",X"3A",X"AE",X"99",X"99",X"99",X"59",X"99",X"99",
		X"F9",X"93",X"93",X"FF",X"FF",X"39",X"33",X"99",X"F9",X"9F",X"7A",X"99",X"FF",X"FA",X"AA",X"99",
		X"F9",X"FA",X"A9",X"9E",X"FF",X"99",X"99",X"9E",X"F9",X"95",X"99",X"9E",X"FF",X"99",X"99",X"9E",
		X"99",X"9A",X"39",X"5E",X"FF",X"9E",X"A9",X"EA",X"99",X"F9",X"A9",X"EE",X"AA",X"EE",X"A9",X"5A",
		X"36",X"EE",X"A9",X"EE",X"A6",X"99",X"A9",X"5E",X"E6",X"EA",X"A9",X"5E",X"E6",X"AE",X"AE",X"E5",
		X"EE",X"AA",X"A3",X"E5",X"9E",X"E9",X"9E",X"9E",X"35",X"AA",X"99",X"99",X"D9",X"D9",X"99",X"FF",
		X"00",X"09",X"99",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"93",X"00",X"00",
		X"99",X"EE",X"00",X"00",X"FF",X"9E",X"99",X"00",X"99",X"F9",X"99",X"00",X"A7",X"9F",X"99",X"00",
		X"AA",X"A9",X"99",X"00",X"AA",X"A7",X"AA",X"00",X"AA",X"AA",X"AA",X"00",X"A9",X"AA",X"A9",X"00",
		X"44",X"AA",X"59",X"00",X"A4",X"AA",X"9A",X"00",X"AA",X"AA",X"9A",X"00",X"AA",X"AA",X"9E",X"00",
		X"A9",X"AA",X"9E",X"00",X"94",X"AA",X"9E",X"00",X"44",X"AA",X"9E",X"00",X"AE",X"AA",X"9E",X"00",
		X"AE",X"AA",X"E5",X"00",X"EE",X"AA",X"AE",X"00",X"EE",X"AA",X"AE",X"00",X"99",X"AE",X"9A",X"00",
		X"FF",X"55",X"59",X"00",X"99",X"99",X"A5",X"00",X"D9",X"F9",X"4A",X"00",X"09",X"99",X"94",X"00",
		X"0D",X"EE",X"99",X"00",X"00",X"E3",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"6E",X"00",X"00",X"00",X"6E",X"00",X"00",X"00",X"6A",X"AE",X"00",X"00",X"3A",X"AA",X"00",X"00",
		X"99",X"A9",X"90",X"00",X"99",X"9A",X"A9",X"50",X"FF",X"A9",X"9E",X"EE",X"99",X"99",X"FA",X"9E",
		X"9F",X"99",X"9F",X"99",X"9F",X"F9",X"A9",X"FA",X"FF",X"F9",X"99",X"9A",X"9F",X"F9",X"A7",X"A9",
		X"9F",X"9A",X"EA",X"99",X"F9",X"9A",X"AE",X"A7",X"F9",X"9A",X"EA",X"EA",X"F9",X"9A",X"AE",X"AE",
		X"99",X"AE",X"EE",X"EA",X"FF",X"AA",X"EE",X"AE",X"FF",X"9A",X"EE",X"EA",X"99",X"99",X"5E",X"AE",
		X"AE",X"99",X"EE",X"AA",X"5E",X"9A",X"E5",X"EA",X"E5",X"9D",X"65",X"AA",X"5E",X"9D",X"AA",X"A7",
		X"EE",X"9D",X"DD",X"5A",X"00",X"EA",X"DD",X"AA",X"00",X"EE",X"DD",X"DD",X"00",X"00",X"AA",X"DD",
		X"00",X"00",X"EE",X"DD",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"95",X"00",X"00",X"00",X"95",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EA",X"00",X"00",X"EA",
		X"E5",X"99",X"9E",X"EE",X"5E",X"EA",X"E9",X"99",X"E5",X"99",X"A9",X"A9",X"AA",X"9A",X"9A",X"9A",
		X"99",X"99",X"A9",X"A9",X"F9",X"99",X"99",X"99",X"F9",X"97",X"A7",X"A7",X"9A",X"95",X"EA",X"AA",
		X"9A",X"A5",X"AE",X"A7",X"9A",X"A5",X"EA",X"AA",X"99",X"E5",X"AE",X"A7",X"99",X"E5",X"EA",X"AA",
		X"9E",X"E5",X"EE",X"A7",X"9E",X"E5",X"EE",X"AA",X"9E",X"A5",X"EE",X"A7",X"9E",X"A5",X"EE",X"AA",
		X"9E",X"95",X"5E",X"A7",X"F9",X"96",X"65",X"5A",X"F9",X"9A",X"AA",X"AA",X"99",X"9D",X"DD",X"DD",
		X"AE",X"9D",X"DD",X"DD",X"5E",X"9D",X"DD",X"DD",X"E5",X"EA",X"AA",X"AA",X"5E",X"EE",X"EE",X"5E",
		X"EE",X"90",X"90",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"F9",X"99",X"00",X"00",X"E9",X"EA",X"00",X"00",
		X"99",X"AA",X"99",X"00",X"99",X"99",X"AA",X"9A",X"99",X"99",X"EE",X"AA",X"99",X"99",X"55",X"99",
		X"99",X"49",X"50",X"55",X"44",X"99",X"99",X"99",X"99",X"93",X"33",X"39",X"AA",X"93",X"EB",X"A3",
		X"AA",X"90",X"3E",X"E9",X"AA",X"90",X"EE",X"99",X"AA",X"00",X"3E",X"09",X"44",X"3F",X"BE",X"99",
		X"E4",X"3F",X"AE",X"99",X"EE",X"9F",X"BE",X"99",X"99",X"95",X"EE",X"99",X"99",X"95",X"BE",X"99",
		X"EE",X"93",X"BB",X"9A",X"EA",X"93",X"99",X"39",X"EE",X"A9",X"55",X"99",X"99",X"99",X"55",X"99",
		X"00",X"EA",X"EE",X"9C",X"00",X"99",X"AE",X"55",X"00",X"00",X"99",X"EE",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"3E",X"00",X"00",X"00",
		X"E3",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A9",
		X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"EE",X"00",X"99",X"AE",X"55",X"00",X"EA",X"EE",X"9C",
		X"99",X"99",X"55",X"99",X"EE",X"A9",X"55",X"99",X"EE",X"93",X"99",X"39",X"EE",X"93",X"BB",X"9A",
		X"99",X"95",X"BE",X"99",X"99",X"95",X"EE",X"99",X"EE",X"9F",X"BE",X"99",X"E4",X"3F",X"AE",X"99",
		X"44",X"3F",X"BE",X"99",X"AA",X"00",X"3E",X"09",X"AA",X"90",X"EE",X"99",X"AA",X"90",X"3E",X"E9",
		X"AA",X"93",X"EB",X"A3",X"99",X"93",X"33",X"39",X"44",X"99",X"99",X"99",X"99",X"49",X"50",X"55",
		X"99",X"99",X"55",X"99",X"99",X"99",X"EE",X"AA",X"99",X"99",X"AA",X"9A",X"99",X"AA",X"99",X"00",
		X"E9",X"EA",X"00",X"00",X"F9",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"40",X"00",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"99",X"90",X"90",X"99",X"99",X"09",X"09",X"22",X"29",X"99",X"99",X"22",X"22",
		X"99",X"99",X"22",X"22",X"33",X"A9",X"22",X"22",X"13",X"39",X"22",X"22",X"A1",X"A9",X"22",X"22",
		X"1A",X"F9",X"22",X"22",X"92",X"22",X"22",X"22",X"23",X"77",X"22",X"22",X"71",X"47",X"22",X"22",
		X"13",X"47",X"22",X"22",X"19",X"46",X"22",X"22",X"19",X"61",X"22",X"22",X"19",X"61",X"22",X"22",
		X"99",X"61",X"22",X"22",X"72",X"61",X"22",X"22",X"11",X"76",X"22",X"22",X"12",X"47",X"22",X"22",
		X"11",X"77",X"22",X"22",X"77",X"47",X"22",X"22",X"23",X"77",X"22",X"22",X"92",X"22",X"22",X"22",
		X"1A",X"F9",X"22",X"22",X"A1",X"29",X"22",X"22",X"13",X"29",X"22",X"22",X"3A",X"A9",X"22",X"22",
		X"99",X"00",X"22",X"22",X"00",X"00",X"22",X"29",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"52",X"00",X"00",X"00",X"11",X"00",X"00",X"55",X"11",X"00",X"00",X"55",X"11",X"00",
		X"00",X"55",X"11",X"50",X"55",X"55",X"11",X"55",X"55",X"55",X"11",X"55",X"55",X"33",X"11",X"33",
		X"55",X"41",X"11",X"33",X"11",X"93",X"39",X"39",X"44",X"33",X"BB",X"41",X"11",X"33",X"99",X"95",
		X"11",X"55",X"99",X"55",X"15",X"55",X"33",X"55",X"55",X"5A",X"51",X"55",X"55",X"5A",X"11",X"55",
		X"FF",X"5A",X"57",X"55",X"FF",X"5A",X"55",X"55",X"1F",X"55",X"55",X"55",X"11",X"55",X"99",X"F5",
		X"11",X"55",X"99",X"95",X"44",X"FF",X"BB",X"11",X"11",X"11",X"FF",X"FF",X"55",X"41",X"11",X"F5",
		X"55",X"55",X"11",X"55",X"F5",X"55",X"11",X"5F",X"F5",X"55",X"11",X"F0",X"00",X"55",X"11",X"00",
		X"00",X"FF",X"11",X"00",X"00",X"FF",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"FF",X"90",X"00",X"00",X"E0",X"F0",X"00",X"00",
		X"33",X"00",X"00",X"00",X"55",X"30",X"00",X"00",X"19",X"95",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",
		X"F9",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"1F",X"50",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E0",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"29",X"00",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"23",X"F3",X"00",X"00",X"22",X"33",X"00",X"00",X"99",X"99",X"99",X"00",
		X"99",X"9F",X"F9",X"00",X"33",X"F3",X"F9",X"00",X"33",X"3F",X"9F",X"00",X"99",X"9F",X"9F",X"00",
		X"92",X"99",X"9F",X"00",X"22",X"F9",X"9F",X"00",X"22",X"F9",X"FF",X"00",X"22",X"99",X"F0",X"00",
		X"29",X"99",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"99",X"90",X"00",X"22",X"99",X"00",X"00",
		X"22",X"99",X"00",X"00",X"22",X"F9",X"00",X"00",X"99",X"99",X"90",X"00",X"22",X"39",X"00",X"00",
		X"22",X"95",X"00",X"00",X"22",X"95",X"00",X"00",X"22",X"95",X"90",X"00",X"22",X"99",X"00",X"00",
		X"11",X"99",X"00",X"00",X"11",X"95",X"90",X"00",X"11",X"95",X"00",X"00",X"11",X"95",X"00",X"00",
		X"11",X"39",X"00",X"00",X"11",X"99",X"90",X"00",X"11",X"F9",X"00",X"00",X"22",X"99",X"00",X"00",
		X"22",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"11",X"99",X"00",X"00",X"11",X"99",X"00",X"00",
		X"11",X"99",X"F0",X"00",X"11",X"F9",X"FF",X"00",X"11",X"F9",X"9F",X"00",X"91",X"99",X"9F",X"00",
		X"99",X"9F",X"9F",X"00",X"33",X"3F",X"9F",X"00",X"33",X"F3",X"F9",X"00",X"99",X"9F",X"F9",X"00",
		X"99",X"99",X"99",X"00",X"22",X"33",X"00",X"00",X"23",X"F3",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"00",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"99",X"00",X"00",X"19",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"99",X"50",X"00",X"00",
		X"F1",X"55",X"00",X"00",X"1F",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"51",X"55",X"00",X"00",
		X"55",X"55",X"00",X"00",X"F5",X"55",X"00",X"00",X"FF",X"15",X"50",X"00",X"FF",X"11",X"55",X"00",
		X"FF",X"11",X"55",X"00",X"FF",X"11",X"55",X"00",X"1F",X"31",X"55",X"00",X"1F",X"53",X"55",X"00",
		X"1F",X"55",X"11",X"00",X"1F",X"99",X"11",X"00",X"11",X"99",X"11",X"00",X"11",X"BB",X"19",X"90",
		X"11",X"99",X"99",X"00",X"11",X"99",X"95",X"00",X"51",X"99",X"12",X"09",X"51",X"99",X"12",X"00",
		X"55",X"99",X"11",X"09",X"55",X"91",X"F1",X"00",X"55",X"B9",X"B1",X"00",X"55",X"BB",X"91",X"00",
		X"55",X"FB",X"99",X"09",X"55",X"FB",X"99",X"00",X"F5",X"1F",X"95",X"09",X"05",X"11",X"5F",X"90",
		X"55",X"35",X"99",X"00",X"95",X"35",X"99",X"90",X"0F",X"33",X"19",X"96",X"00",X"13",X"11",X"96",
		X"00",X"11",X"31",X"00",X"90",X"51",X"31",X"90",X"09",X"F1",X"F3",X"99",X"90",X"FF",X"99",X"99",
		X"00",X"FF",X"FF",X"F6",X"00",X"F9",X"99",X"00",X"00",X"F9",X"9F",X"06",X"00",X"F9",X"FF",X"00",
		X"00",X"F9",X"9F",X"F0",X"00",X"F9",X"3F",X"00",X"00",X"F9",X"3F",X"90",X"00",X"0F",X"13",X"00",
		X"00",X"0F",X"11",X"09",X"00",X"0F",X"F1",X"00",X"00",X"00",X"F2",X"90",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"90",X"00",X"00",X"33",X"99",X"90",X"00",X"15",X"33",X"99",X"00",X"11",X"F3",X"09",X"00",
		X"91",X"5F",X"99",X"00",X"51",X"55",X"33",X"09",X"55",X"5F",X"FF",X"00",X"55",X"15",X"FF",X"99",
		X"55",X"11",X"55",X"99",X"F5",X"11",X"55",X"19",X"FF",X"F1",X"55",X"99",X"FF",X"99",X"11",X"99",
		X"FF",X"95",X"11",X"99",X"1F",X"F5",X"11",X"90",X"11",X"FF",X"11",X"39",X"11",X"FF",X"B1",X"33",
		X"51",X"5F",X"9B",X"F3",X"55",X"FF",X"99",X"5F",X"55",X"FF",X"92",X"5F",X"55",X"FF",X"22",X"55",
		X"F5",X"1F",X"52",X"55",X"FF",X"11",X"55",X"95",X"FF",X"11",X"95",X"19",X"FF",X"11",X"99",X"91",
		X"0F",X"51",X"F9",X"9F",X"00",X"55",X"11",X"9F",X"00",X"F5",X"11",X"FF",X"00",X"55",X"55",X"F8",
		X"00",X"F5",X"55",X"98",X"00",X"FF",X"55",X"11",X"00",X"FF",X"5F",X"51",X"00",X"FF",X"90",X"5F",
		X"55",X"39",X"00",X"00",X"55",X"F9",X"00",X"00",X"55",X"11",X"90",X"00",X"15",X"11",X"00",X"00",
		X"11",X"11",X"09",X"00",X"11",X"19",X"00",X"00",X"F1",X"99",X"00",X"00",X"BB",X"99",X"09",X"00",
		X"BB",X"95",X"00",X"00",X"B9",X"5F",X"09",X"00",X"99",X"15",X"09",X"00",X"99",X"11",X"00",X"00",
		X"99",X"91",X"99",X"00",X"99",X"99",X"F9",X"00",X"B9",X"DF",X"FF",X"00",X"BB",X"DF",X"30",X"90",
		X"1F",X"FF",X"33",X"F0",X"11",X"FF",X"F3",X"00",X"11",X"F9",X"9F",X"00",X"19",X"99",X"91",X"99",
		X"19",X"11",X"8F",X"FF",X"19",X"11",X"F9",X"9F",X"19",X"F9",X"9F",X"F9",X"19",X"F9",X"9F",X"FF",
		X"19",X"F9",X"95",X"3F",X"19",X"F9",X"19",X"39",X"19",X"F9",X"11",X"99",X"19",X"F9",X"FF",X"90",
		X"19",X"FF",X"00",X"90",X"22",X"0F",X"00",X"90",X"00",X"00",X"90",X"09",X"00",X"00",X"99",X"90",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"CC",X"00",X"99",X"00",X"BB",X"99",X"99",X"00",
		X"96",X"99",X"99",X"00",X"9C",X"99",X"99",X"00",X"5A",X"CC",X"99",X"00",X"AA",X"CA",X"99",X"00",
		X"AB",X"E9",X"CC",X"00",X"BE",X"B9",X"EB",X"90",X"EB",X"A9",X"C9",X"99",X"BB",X"A9",X"BE",X"C9",
		X"EE",X"A9",X"EB",X"C9",X"55",X"A9",X"BE",X"49",X"BB",X"A9",X"BB",X"4F",X"BB",X"A9",X"BB",X"44",
		X"BB",X"9B",X"BB",X"59",X"6F",X"9F",X"BB",X"59",X"B6",X"9F",X"BB",X"59",X"9B",X"9F",X"BB",X"59",
		X"C9",X"9F",X"BB",X"59",X"BB",X"9B",X"FB",X"59",X"B6",X"BB",X"BF",X"59",X"BC",X"BB",X"F9",X"54",
		X"9C",X"0B",X"BB",X"40",X"00",X"C0",X"BB",X"40",X"00",X"0C",X"CC",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"90",X"99",X"00",X"09",X"99",X"99",X"00",X"09",X"9C",X"CC",X"00",X"99",X"CA",X"AB",X"40",
		X"0C",X"0A",X"BB",X"40",X"BC",X"AA",X"AB",X"54",X"B6",X"BB",X"BB",X"59",X"BB",X"9B",X"BB",X"59",
		X"C9",X"9B",X"BB",X"59",X"9B",X"9F",X"BB",X"59",X"AA",X"9B",X"BB",X"59",X"AA",X"9F",X"BB",X"59",
		X"BB",X"9B",X"BB",X"59",X"BB",X"A9",X"BB",X"44",X"BB",X"A9",X"BB",X"4F",X"EE",X"A9",X"BE",X"49",
		X"55",X"A9",X"5B",X"C9",X"BB",X"A9",X"B5",X"C9",X"EB",X"B9",X"CF",X"99",X"BE",X"BB",X"EB",X"90",
		X"AF",X"BB",X"CC",X"00",X"BB",X"BB",X"AA",X"00",X"5A",X"CC",X"9A",X"00",X"9C",X"90",X"00",X"00",
		X"96",X"AA",X"00",X"00",X"BB",X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D9",X"00",X"00",X"D9",X"99",X"00",X"09",X"99",X"99",
		X"D9",X"D9",X"99",X"FF",X"35",X"AA",X"99",X"99",X"9E",X"E9",X"9E",X"9E",X"EE",X"AA",X"A3",X"E5",
		X"E6",X"AE",X"AE",X"E5",X"E6",X"EA",X"A9",X"5E",X"A6",X"99",X"A9",X"5E",X"36",X"EE",X"A9",X"EE",
		X"AA",X"EE",X"A9",X"5A",X"99",X"F9",X"A9",X"EE",X"FF",X"9E",X"A9",X"EA",X"99",X"9A",X"39",X"5E",
		X"FF",X"99",X"99",X"9E",X"F9",X"95",X"99",X"9E",X"FF",X"99",X"99",X"9E",X"F9",X"FA",X"A9",X"9E",
		X"FF",X"FA",X"AA",X"99",X"F9",X"9F",X"7A",X"99",X"FF",X"39",X"33",X"99",X"F9",X"93",X"93",X"FF",
		X"99",X"59",X"99",X"99",X"3A",X"AE",X"99",X"99",X"93",X"EA",X"99",X"AA",X"9A",X"AE",X"9A",X"00",
		X"9A",X"A7",X"A0",X"00",X"99",X"AA",X"00",X"00",X"59",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E3",X"99",X"00",X"0D",X"EE",X"99",X"00",
		X"09",X"99",X"94",X"00",X"D9",X"F9",X"4A",X"00",X"99",X"99",X"A5",X"00",X"FF",X"55",X"59",X"00",
		X"99",X"AE",X"9A",X"00",X"EE",X"AA",X"AE",X"00",X"EE",X"AA",X"AE",X"00",X"AE",X"AA",X"E5",X"00",
		X"AE",X"AA",X"9E",X"00",X"44",X"AA",X"9E",X"00",X"94",X"AA",X"9E",X"00",X"A9",X"AA",X"9E",X"00",
		X"AA",X"AA",X"9E",X"00",X"AA",X"AA",X"9A",X"00",X"A4",X"AA",X"9A",X"00",X"44",X"AA",X"59",X"00",
		X"A9",X"AA",X"A9",X"00",X"AA",X"AA",X"AA",X"00",X"AA",X"A7",X"AA",X"00",X"AA",X"A9",X"99",X"00",
		X"A7",X"9F",X"99",X"00",X"99",X"F9",X"99",X"00",X"FF",X"9E",X"99",X"00",X"99",X"EE",X"00",X"00",
		X"99",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"09",X"00",X"00",X"D2",X"99",X"90",X"90",
		X"1D",X"22",X"99",X"99",X"11",X"22",X"22",X"99",X"F1",X"11",X"22",X"22",X"17",X"99",X"22",X"22",
		X"11",X"99",X"99",X"22",X"11",X"99",X"33",X"91",X"EE",X"33",X"11",X"11",X"74",X"33",X"D7",X"91",
		X"74",X"33",X"77",X"99",X"74",X"33",X"77",X"39",X"74",X"33",X"77",X"39",X"75",X"33",X"77",X"39",
		X"7F",X"31",X"77",X"99",X"1D",X"31",X"77",X"99",X"EE",X"91",X"77",X"99",X"11",X"91",X"77",X"99",
		X"11",X"91",X"77",X"99",X"77",X"11",X"57",X"95",X"52",X"99",X"11",X"59",X"22",X"29",X"30",X"99",
		X"99",X"02",X"11",X"99",X"00",X"22",X"22",X"11",X"00",X"00",X"55",X"11",X"00",X"00",X"22",X"11",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"22",X"00",X"00",X"99",X"22",
		X"00",X"99",X"22",X"11",X"00",X"99",X"22",X"11",X"90",X"92",X"22",X"11",X"99",X"02",X"11",X"99",
		X"22",X"29",X"30",X"99",X"44",X"99",X"11",X"99",X"77",X"11",X"77",X"99",X"11",X"91",X"77",X"99",
		X"11",X"91",X"77",X"99",X"EE",X"91",X"77",X"99",X"1D",X"31",X"77",X"99",X"44",X"31",X"77",X"99",
		X"7A",X"33",X"77",X"39",X"A4",X"33",X"77",X"3F",X"74",X"33",X"77",X"F9",X"74",X"33",X"77",X"99",
		X"74",X"FF",X"55",X"91",X"77",X"33",X"11",X"11",X"11",X"99",X"33",X"91",X"11",X"99",X"99",X"22",
		X"17",X"99",X"22",X"52",X"F1",X"11",X"22",X"22",X"11",X"22",X"25",X"00",X"1D",X"22",X"90",X"00",
		X"D2",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"93",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"53",X"00",X"00",
		X"00",X"53",X"00",X"00",X"00",X"53",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"F3",X"00",X"00",
		X"00",X"F3",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"59",X"00",X"00",
		X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"9A",X"90",X"00",X"9B",X"AB",X"A9",X"00",X"9D",X"BD",X"A9",X"00",X"9B",X"BB",X"B9",
		X"00",X"5B",X"5B",X"A9",X"00",X"9A",X"BA",X"B9",X"09",X"D9",X"99",X"EE",X"99",X"EE",X"99",X"99",
		X"DD",X"59",X"E5",X"55",X"99",X"39",X"B9",X"99",X"DD",X"99",X"59",X"E9",X"99",X"99",X"B9",X"9A",
		X"DD",X"99",X"59",X"AB",X"99",X"99",X"B9",X"BA",X"DD",X"99",X"59",X"AB",X"99",X"EE",X"B9",X"BA",
		X"AA",X"BB",X"B9",X"AB",X"AB",X"99",X"B9",X"BA",X"BA",X"99",X"59",X"AB",X"AB",X"99",X"BA",X"9A",
		X"BA",X"99",X"59",X"9A",X"AB",X"99",X"B9",X"F9",X"BA",X"99",X"59",X"99",X"AB",X"B9",X"F5",X"55",
		X"BA",X"5B",X"95",X"55",X"0B",X"A5",X"99",X"55",X"00",X"99",X"99",X"99",X"00",X"9A",X"BA",X"9B",
		X"00",X"AB",X"AB",X"9A",X"00",X"9B",X"BB",X"9B",X"00",X"B5",X"B5",X"9A",X"00",X"9B",X"AB",X"90",
		X"99",X"99",X"00",X"00",X"AB",X"AB",X"00",X"00",X"9D",X"BD",X"90",X"00",X"9B",X"BB",X"90",X"00",
		X"5B",X"5B",X"90",X"00",X"9A",X"BA",X"90",X"00",X"DD",X"DD",X"90",X"00",X"ED",X"DD",X"90",X"00",
		X"EB",X"BB",X"90",X"00",X"ED",X"DD",X"90",X"00",X"EB",X"BB",X"90",X"00",X"ED",X"DD",X"90",X"00",
		X"EB",X"BB",X"90",X"00",X"EB",X"DB",X"90",X"00",X"EB",X"BB",X"90",X"00",X"EB",X"BB",X"90",X"00",
		X"EB",X"BA",X"90",X"00",X"EB",X"BB",X"90",X"00",X"EB",X"AB",X"90",X"00",X"EB",X"BB",X"90",X"00",
		X"EA",X"AA",X"90",X"00",X"EB",X"BB",X"90",X"00",X"EA",X"AA",X"90",X"00",X"E9",X"B9",X"90",X"00",
		X"EA",X"C5",X"90",X"00",X"59",X"B9",X"90",X"00",X"99",X"99",X"90",X"00",X"9B",X"AB",X"90",X"00",
		X"9A",X"BA",X"A0",X"00",X"9B",X"BB",X"A0",X"00",X"B5",X"B5",X"00",X"00",X"AB",X"AB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"FF",X"BB",X"BB",X"00",X"FF",X"BB",X"BB",X"00",
		X"FF",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"BB",X"00",X"BB",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BF",X"00",
		X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BF",X"00",X"BB",X"0B",X"BF",X"00",
		X"BB",X"0B",X"BF",X"00",X"BB",X"0B",X"BF",X"00",X"BB",X"0B",X"BF",X"00",X"FB",X"BB",X"BF",X"00",
		X"FF",X"BB",X"BF",X"00",X"BF",X"BB",X"BF",X"00",X"BB",X"BB",X"BF",X"00",X"0B",X"FB",X"FF",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",
		X"BB",X"FF",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"B0",X"FB",X"00",X"BB",X"00",X"BB",X"00",
		X"FF",X"00",X"0B",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"0B",X"00",X"00",
		X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"FB",X"00",
		X"BB",X"BB",X"BF",X"00",X"BB",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"BB",X"00",X"BB",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"B0",X"00",X"BF",X"00",X"FB",X"00",
		X"BB",X"0B",X"BF",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",
		X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",
		X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"BF",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"0B",X"BB",X"FF",X"00",
		X"BB",X"BB",X"BF",X"00",X"FB",X"BB",X"BB",X"00",X"BB",X"B0",X"BB",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"00",X"0B",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"FB",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"0B",X"00",X"00",
		X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"FB",X"00",X"BB",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"BB",X"00",X"BB",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"FB",X"0F",X"BB",X"00",X"FB",X"0F",X"BF",X"00",
		X"FF",X"0F",X"BB",X"00",X"FF",X"0F",X"BB",X"00",X"BF",X"0B",X"FF",X"00",X"FB",X"0B",X"FF",X"00",
		X"BF",X"0B",X"FF",X"00",X"BF",X"0B",X"BF",X"00",X"BF",X"0B",X"BF",X"00",X"BB",X"BB",X"BF",X"00",
		X"BB",X"BF",X"BF",X"00",X"BB",X"BB",X"BF",X"00",X"BB",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FB",X"B0",X"00",X"00",X"FF",X"BB",X"00",X"0B",X"BB",X"BB",X"00",
		X"BB",X"BB",X"FB",X"00",X"BB",X"BB",X"BF",X"00",X"FF",X"B0",X"BB",X"00",X"FB",X"00",X"BB",X"00",
		X"BB",X"00",X"0B",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"FB",X"BB",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"BF",X"00",X"00",X"FB",X"0B",X"00",X"00",
		X"FB",X"0B",X"00",X"00",X"FB",X"0B",X"00",X"00",X"FF",X"0B",X"00",X"00",X"BF",X"0B",X"00",X"00",
		X"FB",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"FF",X"BB",X"BB",X"00",X"FF",X"BB",X"BB",X"00",
		X"FF",X"FB",X"BB",X"00",X"BB",X"FF",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"FF",X"00",
		X"BB",X"00",X"BB",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"B0",X"00",X"BB",X"00",X"BB",X"00",
		X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"FF",X"00",
		X"BB",X"0B",X"FB",X"00",X"BB",X"0B",X"BF",X"00",X"BB",X"0B",X"BF",X"00",X"FB",X"0B",X"BF",X"00",
		X"FB",X"0B",X"BF",X"00",X"FB",X"0B",X"BF",X"00",X"FB",X"0B",X"BF",X"00",X"FF",X"BB",X"BF",X"00",
		X"FF",X"BB",X"BF",X"00",X"FF",X"BB",X"BF",X"00",X"FF",X"BB",X"BF",X"00",X"0B",X"FB",X"FF",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"0B",X"FF",X"BB",X"00",
		X"BB",X"FF",X"BB",X"00",X"BB",X"FB",X"BB",X"00",X"BB",X"B0",X"FF",X"00",X"BB",X"00",X"BB",X"00",
		X"FF",X"00",X"0B",X"00",X"FF",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"0B",X"00",X"00",
		X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"FB",X"0B",X"00",X"00",X"FB",X"0B",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",X"00",
		X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",X"00",X"00",
		X"11",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"01",X"00",
		X"00",X"11",X"01",X"00",X"00",X"11",X"01",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"10",X"00",
		X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"01",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"11",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"11",X"11",X"01",X"00",X"11",X"11",X"01",X"00",X"00",X"11",X"01",X"00",X"00",X"11",X"01",X"00",
		X"00",X"11",X"01",X"00",X"00",X"11",X"01",X"00",X"00",X"11",X"01",X"00",X"00",X"11",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"0E",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"02",X"A0",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"09",X"A0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"09",X"AA",X"00",X"00",X"05",X"0A",X"00",X"00",X"25",X"0A",X"00",
		X"00",X"22",X"00",X"00",X"00",X"02",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"25",X"A0",X"00",
		X"00",X"22",X"AA",X"00",X"00",X"02",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",
		X"00",X"0E",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"02",X"A0",X"00",X"00",X"22",X"00",X"00",
		X"00",X"22",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"09",X"AA",X"00",X"00",X"EE",X"AA",X"00",
		X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"05",X"9F",X"00",X"00",X"0F",X"99",X"00",X"00",X"B9",X"99",X"00",
		X"00",X"59",X"99",X"00",X"00",X"5B",X"99",X"00",X"00",X"0B",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"09",X"09",X"99",X"09",X"99",X"99",X"90",
		X"55",X"99",X"99",X"59",X"EE",X"EE",X"EE",X"EE",X"BB",X"BB",X"BB",X"BB",X"44",X"5F",X"99",X"55",
		X"77",X"95",X"9F",X"FE",X"45",X"99",X"FF",X"59",X"55",X"99",X"FF",X"95",X"FF",X"99",X"FF",X"B5",
		X"E5",X"99",X"FF",X"55",X"EE",X"39",X"FF",X"95",X"F5",X"39",X"FF",X"95",X"F5",X"39",X"FF",X"95",
		X"F5",X"39",X"FF",X"95",X"FF",X"39",X"FF",X"95",X"FF",X"39",X"FF",X"95",X"FF",X"39",X"FF",X"55",
		X"F5",X"39",X"FF",X"35",X"55",X"33",X"FF",X"95",X"55",X"93",X"FF",X"59",X"77",X"95",X"9F",X"55",
		X"44",X"5F",X"99",X"55",X"BF",X"BB",X"BB",X"BB",X"FF",X"FF",X"FF",X"FF",X"55",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"F9",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"F5",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
