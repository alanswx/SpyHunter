library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_sp_bits_2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_sp_bits_2 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"22",X"20",X"00",X"00",X"22",X"10",X"00",X"00",X"22",X"10",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"20",X"00",X"00",X"02",X"20",X"00",X"00",X"22",X"20",
		X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",
		X"00",X"00",X"99",X"90",X"00",X"AA",X"AA",X"EA",X"00",X"EB",X"AA",X"BE",X"00",X"BB",X"AA",X"EB",
		X"00",X"99",X"99",X"BE",X"9B",X"AA",X"99",X"EE",X"0E",X"AA",X"BB",X"BB",X"0B",X"A9",X"BB",X"BB",
		X"BB",X"A9",X"5B",X"5B",X"BB",X"AA",X"55",X"55",X"BB",X"A9",X"FA",X"55",X"BB",X"55",X"AA",X"F5",
		X"BB",X"A9",X"FA",X"55",X"BB",X"A9",X"55",X"55",X"BB",X"AF",X"5B",X"5B",X"0B",X"F9",X"BB",X"BB",
		X"0C",X"AA",X"BB",X"BB",X"9B",X"AA",X"A9",X"EB",X"00",X"99",X"9A",X"BE",X"00",X"BB",X"9A",X"EB",
		X"00",X"EB",X"AA",X"BE",X"00",X"AA",X"AA",X"EA",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",X"EB",X"AA",X"00",X"00",
		X"BE",X"EB",X"AA",X"00",X"BB",X"B5",X"EE",X"AA",X"55",X"55",X"B6",X"B5",X"5F",X"FF",X"FF",X"55",
		X"55",X"55",X"B5",X"B6",X"BB",X"B5",X"EE",X"AA",X"BE",X"EB",X"AA",X"00",X"EB",X"AA",X"00",X"00",
		X"BE",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"0A",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",X"A9",X"90",
		X"00",X"A9",X"BA",X"99",X"00",X"AA",X"BA",X"99",X"00",X"AA",X"BA",X"00",X"00",X"AA",X"BA",X"00",
		X"99",X"A9",X"BA",X"00",X"99",X"59",X"EE",X"99",X"00",X"5B",X"BB",X"99",X"00",X"BB",X"BB",X"9E",
		X"00",X"BB",X"5B",X"BE",X"00",X"BB",X"55",X"EB",X"00",X"BB",X"A5",X"BE",X"00",X"9B",X"AF",X"BB",
		X"00",X"9B",X"6F",X"BB",X"00",X"99",X"55",X"BB",X"00",X"B9",X"55",X"5B",X"00",X"BB",X"BB",X"55",
		X"00",X"BB",X"BB",X"F5",X"00",X"AB",X"AB",X"FF",X"00",X"A9",X"AA",X"5F",X"00",X"90",X"A9",X"55",
		X"00",X"99",X"99",X"BB",X"00",X"99",X"99",X"BB",X"00",X"99",X"99",X"EB",X"00",X"09",X"09",X"BE",
		X"00",X"00",X"00",X"EB",X"00",X"00",X"90",X"AA",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"5B",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"5F",X"A0",X"00",X"00",X"BB",X"BA",X"00",X"00",X"AA",X"BB",X"00",X"00",
		X"AA",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"AB",X"A0",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"A9",X"00",X"00",X"BB",X"AA",X"09",X"00",X"BB",X"AA",X"99",X"00",
		X"BB",X"A9",X"90",X"00",X"BA",X"AA",X"90",X"00",X"BA",X"A9",X"90",X"00",X"BA",X"99",X"99",X"00",
		X"AA",X"BB",X"A9",X"00",X"9F",X"5B",X"A9",X"00",X"B9",X"55",X"A9",X"00",X"B9",X"5F",X"AA",X"00",
		X"BB",X"FF",X"AA",X"90",X"BB",X"FF",X"AA",X"90",X"BB",X"5A",X"AA",X"99",X"BB",X"5A",X"9A",X"99",
		X"AB",X"55",X"99",X"09",X"AB",X"55",X"99",X"00",X"09",X"B5",X"B9",X"00",X"99",X"BB",X"BB",X"00",
		X"00",X"BB",X"BE",X"00",X"00",X"BB",X"BB",X"00",X"00",X"9B",X"BE",X"00",X"90",X"9B",X"BB",X"00",
		X"90",X"99",X"BB",X"00",X"99",X"9B",X"5B",X"00",X"09",X"BE",X"5B",X"00",X"09",X"AB",X"5B",X"00",
		X"00",X"AA",X"F5",X"00",X"00",X"0A",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"B5",X"00",
		X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",
		X"00",X"00",X"00",X"BC",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"BB",X"00",X"00",X"BC",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"AB",X"00",X"00",X"BB",X"AA",X"00",X"00",X"BA",X"AA",X"00",
		X"00",X"BF",X"AA",X"00",X"00",X"AF",X"AA",X"00",X"00",X"AA",X"AA",X"00",X"00",X"AA",X"99",X"00",
		X"00",X"99",X"BB",X"00",X"00",X"99",X"BB",X"00",X"00",X"9B",X"5B",X"00",X"00",X"BB",X"55",X"00",
		X"00",X"BB",X"5B",X"99",X"00",X"9B",X"55",X"90",X"00",X"99",X"55",X"00",X"00",X"99",X"5B",X"00",
		X"00",X"99",X"55",X"00",X"00",X"99",X"5B",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"00",
		X"00",X"99",X"5B",X"00",X"00",X"99",X"55",X"00",X"00",X"99",X"55",X"99",X"00",X"BB",X"5B",X"99",
		X"00",X"EB",X"55",X"09",X"00",X"BE",X"5B",X"00",X"00",X"EB",X"BB",X"00",X"00",X"BE",X"5B",X"00",
		X"00",X"EB",X"BB",X"00",X"00",X"BE",X"BB",X"00",X"00",X"AB",X"BB",X"00",X"00",X"AE",X"BE",X"00",
		X"00",X"0A",X"BB",X"00",X"00",X"0A",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BE",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",X"00",
		X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",X"00",
		X"00",X"00",X"EA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"50",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"05",X"00",X"55",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",
		X"00",X"35",X"35",X"00",X"00",X"05",X"03",X"00",X"00",X"05",X"05",X"F0",X"00",X"05",X"05",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F5",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"05",X"F0",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"FF",X"F5",X"00",X"00",X"F5",X"F0",X"00",X"00",X"5F",X"53",X"00",
		X"00",X"50",X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"05",X"3F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"05",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"0F",X"90",X"00",X"90",
		X"05",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"55",X"09",X"90",X"00",X"95",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"00",X"00",X"00",
		X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"F1",X"1F",X"00",X"00",X"16",X"FF",
		X"00",X"00",X"04",X"01",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"31",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"91",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FA",X"A0",X"00",
		X"00",X"FA",X"A0",X"00",X"00",X"5A",X"A0",X"00",X"05",X"5A",X"00",X"00",X"0F",X"5A",X"0F",X"00",
		X"0F",X"AA",X"F5",X"00",X"0F",X"5A",X"F5",X"00",X"00",X"5A",X"F5",X"00",X"00",X"5A",X"55",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"F5",X"55",X"00",X"00",X"F5",X"55",X"00",X"00",X"F5",X"55",X"00",X"00",X"55",X"F5",X"00",
		X"00",X"0F",X"5F",X"00",X"00",X"0F",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"5F",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",X"99",X"00",
		X"09",X"00",X"99",X"00",X"99",X"09",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"09",X"99",X"00",
		X"99",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"90",X"00",
		X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"D9",X"99",X"99",X"00",X"99",X"99",X"D9",X"00",X"99",X"99",X"D9",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"9D",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"35",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"03",X"E3",X"00",X"00",X"55",X"E3",X"00",X"00",X"F5",X"33",X"00",
		X"35",X"F5",X"55",X"00",X"55",X"F5",X"55",X"00",X"F0",X"FF",X"EE",X"00",X"FF",X"50",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"30",X"55",X"30",X"35",X"03",X"55",X"30",X"55",X"5E",X"F5",X"00",
		X"F0",X"5E",X"F5",X"00",X"00",X"E5",X"FF",X"00",X"00",X"55",X"EF",X"00",X"00",X"55",X"EF",X"00",
		X"00",X"0F",X"EE",X"00",X"00",X"0F",X"30",X"00",X"00",X"0F",X"33",X"00",X"00",X"00",X"53",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"30",X"30",X"00",X"55",X"E3",X"30",
		X"00",X"55",X"5E",X"E3",X"00",X"55",X"5E",X"5E",X"00",X"F5",X"5E",X"55",X"00",X"55",X"55",X"55",
		X"00",X"5F",X"55",X"55",X"00",X"F5",X"5F",X"50",X"00",X"5F",X"E5",X"30",X"00",X"55",X"55",X"33",
		X"00",X"F5",X"55",X"EE",X"00",X"F5",X"5E",X"05",X"00",X"05",X"55",X"55",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"5F",X"55",X"00",X"E5",X"55",X"55",X"00",X"5E",X"5F",X"00",
		X"00",X"5E",X"F5",X"00",X"00",X"55",X"FF",X"00",X"00",X"E5",X"3F",X"30",X"00",X"55",X"00",X"E3",
		X"00",X"55",X"00",X"33",X"00",X"F5",X"30",X"53",X"00",X"55",X"30",X"00",X"00",X"F5",X"30",X"00",
		X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"09",X"00",X"00",X"EE",X"00",X"00",X"00",X"BB",X"99",X"00",X"00",X"44",X"99",X"00",
		X"05",X"77",X"99",X"90",X"59",X"55",X"EE",X"90",X"59",X"55",X"BB",X"99",X"5F",X"FF",X"F9",X"E0",
		X"5F",X"B5",X"59",X"BE",X"5F",X"5E",X"55",X"FB",X"5F",X"55",X"9F",X"FB",X"FF",X"5B",X"FF",X"51",
		X"F5",X"55",X"FF",X"99",X"F5",X"55",X"FF",X"99",X"55",X"55",X"FF",X"55",X"F5",X"F5",X"FF",X"FF",
		X"F3",X"5F",X"FF",X"F5",X"FF",X"55",X"FF",X"59",X"FF",X"59",X"FF",X"99",X"B4",X"55",X"FF",X"99",
		X"EF",X"55",X"FF",X"99",X"0F",X"77",X"FF",X"99",X"00",X"45",X"FF",X"99",X"00",X"BB",X"55",X"99",
		X"00",X"FF",X"99",X"99",X"00",X"00",X"99",X"59",X"00",X"00",X"B9",X"55",X"00",X"00",X"FB",X"95",
		X"00",X"00",X"0F",X"55",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"EA",X"90",X"00",X"00",X"5E",X"00",X"00",X"00",
		X"5E",X"90",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"90",X"00",X"00",X"55",X"00",X"00",X"00",
		X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",
		X"E5",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",
		X"A5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"19",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F2",X"00",X"00",X"00",X"FF",X"90",X"00",
		X"00",X"33",X"09",X"00",X"00",X"3F",X"99",X"00",X"00",X"5F",X"99",X"00",X"02",X"5F",X"99",X"00",
		X"22",X"95",X"A9",X"00",X"2F",X"B5",X"A9",X"00",X"2F",X"B5",X"EA",X"00",X"25",X"BB",X"EA",X"00",
		X"E7",X"5B",X"EA",X"00",X"E7",X"55",X"EE",X"00",X"A4",X"5B",X"4E",X"00",X"A4",X"55",X"4E",X"00",
		X"AE",X"55",X"4E",X"00",X"AE",X"55",X"43",X"00",X"AA",X"55",X"53",X"00",X"0A",X"55",X"53",X"00",
		X"0A",X"59",X"F3",X"00",X"0A",X"99",X"F9",X"00",X"00",X"99",X"F9",X"00",X"00",X"99",X"59",X"00",
		X"00",X"99",X"F9",X"00",X"00",X"99",X"F9",X"00",X"00",X"95",X"F5",X"90",X"00",X"9F",X"FF",X"90",
		X"00",X"5F",X"FF",X"99",X"00",X"9F",X"FF",X"99",X"00",X"9F",X"FF",X"99",X"00",X"95",X"FF",X"99",
		X"00",X"99",X"FF",X"99",X"00",X"99",X"FF",X"A9",X"00",X"99",X"99",X"A9",X"00",X"99",X"99",X"AA",
		X"00",X"E5",X"99",X"EA",X"00",X"E5",X"99",X"EA",X"00",X"E7",X"99",X"4A",X"00",X"E7",X"99",X"44",
		X"00",X"EE",X"99",X"4A",X"00",X"AE",X"99",X"3A",X"00",X"AE",X"99",X"3A",X"00",X"AE",X"99",X"AA",
		X"00",X"0A",X"33",X"AA",X"00",X"0A",X"55",X"11",X"00",X"00",X"55",X"19",X"00",X"00",X"55",X"19",
		X"00",X"00",X"44",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"15",X"90",X"00",X"00",X"15",X"90",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"BB",X"00",X"0F",X"00",X"5B",X"00",X"0F",X"00",X"5B",X"00",X"0F",X"B0",X"B0",
		X"00",X"0F",X"5B",X"BB",X"00",X"5F",X"E0",X"5B",X"00",X"5F",X"B0",X"50",X"00",X"F5",X"00",X"B0",
		X"00",X"05",X"00",X"B0",X"00",X"05",X"B0",X"00",X"00",X"5B",X"B0",X"00",X"00",X"5B",X"B0",X"00",
		X"00",X"5F",X"5B",X"00",X"00",X"F5",X"5B",X"00",X"00",X"55",X"BB",X"00",X"00",X"55",X"BB",X"00",
		X"00",X"55",X"5B",X"00",X"00",X"FF",X"F5",X"00",X"00",X"55",X"5B",X"00",X"00",X"5B",X"BB",X"00",
		X"00",X"BB",X"BE",X"00",X"00",X"BB",X"BB",X"00",X"00",X"F5",X"5B",X"00",X"00",X"0F",X"05",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"55",X"50",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"B5",X"55",X"00",X"00",X"5B",X"BB",X"00",X"00",X"55",X"BB",X"00",X"00",X"55",X"B5",X"00",
		X"00",X"55",X"5F",X"00",X"00",X"F5",X"B5",X"00",X"00",X"FF",X"5F",X"00",X"00",X"55",X"B5",X"00",
		X"00",X"05",X"55",X"00",X"00",X"05",X"B5",X"00",X"00",X"05",X"BB",X"00",X"0F",X"05",X"BB",X"00",
		X"05",X"00",X"55",X"00",X"0F",X"00",X"B0",X"00",X"0F",X"0F",X"B0",X"00",X"0F",X"05",X"B0",X"00",
		X"00",X"05",X"B0",X"00",X"00",X"05",X"00",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"99",X"99",X"00",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"A9",X"AA",X"99",X"90",X"A9",X"EE",X"9E",X"00",X"AA",X"55",X"99",X"09",
		X"7A",X"55",X"99",X"99",X"74",X"55",X"FF",X"99",X"57",X"55",X"FF",X"A5",X"F7",X"59",X"FF",X"99",
		X"A5",X"55",X"FF",X"55",X"AA",X"95",X"FF",X"95",X"9A",X"33",X"F9",X"95",X"AA",X"33",X"F9",X"95",
		X"A5",X"33",X"99",X"95",X"A5",X"33",X"9F",X"95",X"55",X"33",X"9F",X"95",X"55",X"33",X"9F",X"55",
		X"FF",X"33",X"9A",X"99",X"57",X"93",X"00",X"55",X"34",X"99",X"00",X"99",X"AA",X"79",X"33",X"99",
		X"A3",X"0A",X"33",X"F4",X"A3",X"0A",X"93",X"EE",X"00",X"0A",X"F9",X"AA",X"09",X"00",X"FF",X"99",
		X"09",X"00",X"9F",X"99",X"09",X"00",X"FF",X"09",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",X"09",X"09",X"00",X"99",X"99",X"99",
		X"09",X"55",X"99",X"5F",X"EE",X"EE",X"EE",X"EE",X"EB",X"BB",X"BB",X"BB",X"E4",X"42",X"99",X"11",
		X"F7",X"77",X"99",X"99",X"F3",X"55",X"55",X"99",X"F5",X"55",X"FF",X"55",X"55",X"55",X"FF",X"F5",
		X"F5",X"55",X"FF",X"59",X"F5",X"B5",X"FF",X"59",X"F5",X"55",X"FF",X"59",X"F5",X"55",X"FF",X"59",
		X"F5",X"55",X"FF",X"59",X"F5",X"55",X"FF",X"59",X"F5",X"FF",X"FF",X"59",X"F5",X"55",X"FF",X"59",
		X"55",X"55",X"FF",X"F5",X"F5",X"55",X"FF",X"55",X"F3",X"55",X"55",X"99",X"FF",X"77",X"99",X"99",
		X"FF",X"42",X"99",X"11",X"EF",X"BB",X"BB",X"BB",X"EE",X"FF",X"FF",X"FF",X"00",X"55",X"00",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"BB",X"90",X"00",X"00",
		X"44",X"09",X"00",X"00",X"E3",X"99",X"00",X"00",X"5E",X"90",X"00",X"00",X"5B",X"99",X"00",X"00",
		X"B5",X"90",X"00",X"00",X"5B",X"99",X"00",X"00",X"B5",X"90",X"00",X"00",X"55",X"99",X"00",X"00",
		X"55",X"90",X"00",X"00",X"55",X"99",X"00",X"00",X"55",X"90",X"00",X"00",X"55",X"09",X"00",X"00",
		X"55",X"90",X"00",X"00",X"F4",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"0C",X"99",X"C9",X"CC",X"C9",X"EB",X"0C",X"BB",X"65",X"CA",X"BE",X"9B",X"65",X"AA",X"AA",X"C9",
		X"65",X"BE",X"EB",X"BC",X"99",X"EB",X"BE",X"B9",X"5A",X"EB",X"BB",X"BB",X"5E",X"BB",X"BB",X"9B",
		X"5E",X"BB",X"BB",X"9A",X"FE",X"EE",X"B5",X"9A",X"F5",X"5F",X"BB",X"9A",X"FE",X"BB",X"5B",X"9A",
		X"5E",X"BB",X"B5",X"99",X"FE",X"BB",X"5B",X"9B",X"5E",X"BB",X"BF",X"BB",X"99",X"BB",X"FB",X"B9",
		X"65",X"96",X"BB",X"BC",X"65",X"BB",X"6F",X"CB",X"65",X"CC",X"BB",X"9B",X"CB",X"BB",X"0C",X"BB",
		X"0C",X"99",X"C9",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"77",X"99",X"99",X"00",X"77",X"DD",X"99",
		X"00",X"76",X"AD",X"99",X"00",X"07",X"DA",X"99",X"00",X"97",X"DD",X"99",X"04",X"19",X"AD",X"94",
		X"E6",X"11",X"7A",X"95",X"96",X"11",X"7A",X"55",X"E6",X"F1",X"7A",X"55",X"96",X"11",X"7A",X"95",
		X"04",X"17",X"7D",X"04",X"00",X"07",X"DD",X"00",X"00",X"97",X"DA",X"00",X"00",X"77",X"AD",X"00",
		X"00",X"76",X"D7",X"00",X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"7A",X"AA",X"AA",
		X"00",X"AE",X"99",X"99",X"0F",X"EE",X"A9",X"99",X"0F",X"9E",X"99",X"99",X"0F",X"9E",X"99",X"A3",
		X"0F",X"9E",X"9A",X"33",X"0F",X"95",X"53",X"FF",X"0F",X"99",X"7A",X"F5",X"0F",X"F9",X"AA",X"55",
		X"0F",X"F3",X"AA",X"55",X"0F",X"FA",X"AA",X"55",X"0F",X"F9",X"99",X"55",X"0F",X"FF",X"55",X"50",
		X"0F",X"FE",X"AA",X"FF",X"0F",X"FE",X"AA",X"F5",X"0F",X"FE",X"EA",X"55",X"0F",X"F9",X"AE",X"55",
		X"0F",X"99",X"EA",X"F5",X"0F",X"AA",X"5E",X"FF",X"0F",X"9E",X"9E",X"FF",X"0F",X"95",X"99",X"A3",
		X"0F",X"9E",X"99",X"EE",X"0F",X"EE",X"A9",X"99",X"00",X"EE",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"F5",X"D9",X"D9",X"00",X"D9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"99",X"99",X"39",X"0F",
		X"99",X"9A",X"E3",X"0F",X"99",X"99",X"99",X"90",X"F9",X"F9",X"99",X"90",X"99",X"99",X"99",X"40",
		X"0A",X"77",X"59",X"90",X"AA",X"AA",X"75",X"90",X"AA",X"AA",X"A7",X"50",X"AA",X"99",X"A5",X"90",
		X"AA",X"44",X"A7",X"90",X"AA",X"49",X"A7",X"90",X"AA",X"9A",X"AA",X"90",X"AA",X"94",X"AA",X"90",
		X"AA",X"49",X"AA",X"90",X"AA",X"94",X"AA",X"90",X"EA",X"9A",X"AE",X"90",X"AA",X"49",X"A5",X"90",
		X"EA",X"44",X"AE",X"90",X"AE",X"AE",X"E5",X"50",X"EE",X"EA",X"E5",X"90",X"EE",X"EE",X"59",X"90",
		X"99",X"99",X"99",X"40",X"F9",X"F9",X"99",X"90",X"99",X"99",X"99",X"90",X"99",X"9A",X"E3",X"0F",
		X"D9",X"D9",X"39",X"0F",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"E9",
		X"09",X"EE",X"AE",X"AA",X"09",X"EA",X"9E",X"E3",X"09",X"EA",X"39",X"53",X"99",X"99",X"53",X"33",
		X"94",X"99",X"F0",X"99",X"99",X"99",X"5F",X"3B",X"55",X"44",X"55",X"EE",X"99",X"4A",X"FF",X"EA",
		X"55",X"91",X"FF",X"EE",X"99",X"94",X"FF",X"AE",X"55",X"49",X"FF",X"EE",X"99",X"94",X"FF",X"EA",
		X"55",X"91",X"F5",X"EE",X"99",X"49",X"55",X"EE",X"55",X"44",X"55",X"EE",X"99",X"EE",X"5F",X"BB",
		X"94",X"99",X"F5",X"99",X"99",X"99",X"53",X"33",X"09",X"A9",X"39",X"53",X"09",X"AA",X"9E",X"E3",
		X"09",X"EE",X"AE",X"AA",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"90",X"90",X"99",X"00",X"09",X"02",X"92",X"09",X"99",X"99",X"22",
		X"99",X"99",X"99",X"22",X"21",X"A3",X"99",X"22",X"17",X"33",X"99",X"22",X"17",X"AA",X"29",X"22",
		X"31",X"3F",X"29",X"22",X"29",X"99",X"29",X"22",X"33",X"52",X"29",X"22",X"29",X"52",X"29",X"22",
		X"97",X"52",X"29",X"22",X"97",X"22",X"29",X"22",X"97",X"27",X"29",X"22",X"97",X"27",X"29",X"22",
		X"99",X"27",X"29",X"22",X"97",X"27",X"29",X"22",X"97",X"27",X"29",X"22",X"97",X"22",X"29",X"22",
		X"97",X"F2",X"29",X"22",X"29",X"F2",X"29",X"22",X"33",X"F9",X"29",X"22",X"39",X"92",X"29",X"22",
		X"21",X"3F",X"29",X"22",X"17",X"AA",X"29",X"22",X"17",X"33",X"09",X"22",X"21",X"A3",X"09",X"22",
		X"99",X"00",X"09",X"22",X"00",X"00",X"02",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"99",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"39",X"33",X"30",X"00",
		X"39",X"93",X"90",X"00",X"30",X"03",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"03",X"00",X"00",
		X"39",X"03",X"00",X"00",X"33",X"33",X"30",X"00",X"99",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"90",X"00",X"33",X"33",X"30",X"00",X"39",X"03",X"00",X"00",
		X"39",X"03",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"03",X"00",X"00",X"39",X"93",X"90",X"00",
		X"39",X"93",X"30",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",
		X"00",X"99",X"09",X"99",X"09",X"99",X"92",X"22",X"92",X"22",X"22",X"22",X"2D",X"22",X"22",X"22",
		X"F2",X"11",X"99",X"99",X"67",X"11",X"33",X"39",X"27",X"19",X"11",X"11",X"21",X"19",X"D7",X"A0",
		X"21",X"19",X"77",X"D1",X"21",X"19",X"77",X"D1",X"21",X"19",X"77",X"71",X"21",X"19",X"77",X"51",
		X"21",X"19",X"77",X"71",X"21",X"19",X"77",X"71",X"21",X"59",X"57",X"51",X"21",X"19",X"77",X"71",
		X"2D",X"1F",X"57",X"51",X"2E",X"19",X"F7",X"71",X"27",X"19",X"11",X"11",X"67",X"11",X"33",X"39",
		X"F2",X"77",X"99",X"99",X"22",X"22",X"22",X"22",X"90",X"22",X"25",X"55",X"00",X"99",X"02",X"22",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"17",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"71",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"F1",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"09",X"09",X"90",X"99",
		X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"09",X"99",X"99",X"09",
		X"09",X"09",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"05",X"55",X"30",X"55",X"55",X"55",X"E3",X"55",
		X"55",X"55",X"5E",X"E5",X"55",X"55",X"5E",X"5E",X"55",X"F5",X"5E",X"55",X"5F",X"55",X"55",X"55",
		X"55",X"5F",X"55",X"55",X"F5",X"F5",X"5F",X"55",X"F5",X"5F",X"E5",X"55",X"5F",X"55",X"55",X"55",
		X"5F",X"F5",X"55",X"E5",X"55",X"F5",X"55",X"55",X"5F",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",
		X"5F",X"55",X"55",X"55",X"55",X"55",X"5F",X"55",X"55",X"E5",X"55",X"55",X"F5",X"5E",X"5F",X"55",
		X"55",X"5E",X"F5",X"55",X"F5",X"55",X"FF",X"55",X"F5",X"E5",X"5F",X"55",X"5F",X"55",X"55",X"E5",
		X"5F",X"55",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",X"55",X"55",X"F5",X"55",X"55",
		X"55",X"55",X"35",X"55",X"55",X"F5",X"00",X"55",X"55",X"0F",X"00",X"00",X"55",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"39",X"00",X"00",X"0F",X"99",X"00",X"00",X"93",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"90",
		X"00",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"90",X"90",X"00",
		X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",
		X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",
		X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",
		X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",
		X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"91",X"00",X"00",X"19",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"01",X"19",X"00",X"00",X"00",X"19",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"D0",X"00",
		X"00",X"00",X"D0",X"00",X"00",X"09",X"D9",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"91",X"00",
		X"00",X"11",X"01",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"11",X"11",X"00",X"00",X"F1",X"10",X"00",X"99",X"FD",X"00",X"00",X"F9",X"9D",X"00",
		X"00",X"FF",X"9D",X"20",X"00",X"00",X"D0",X"00",X"99",X"00",X"60",X"11",X"11",X"10",X"0F",X"11",
		X"11",X"10",X"9F",X"11",X"00",X"11",X"F0",X"19",X"00",X"01",X"00",X"99",X"00",X"91",X"11",X"90",
		X"00",X"91",X"11",X"02",X"00",X"91",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"10",X"11",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"22",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"10",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"60",X"00",X"99",X"11",X"06",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"66",X"00",X"00",X"44",X"40",X"00",X"0F",X"44",X"11",X"66",X"00",
		X"04",X"11",X"00",X"90",X"00",X"11",X"00",X"96",X"00",X"44",X"66",X"00",X"00",X"41",X"66",X"60",
		X"00",X"11",X"00",X"06",X"00",X"40",X"00",X"00",X"00",X"11",X"00",X"60",X"00",X"44",X"16",X"06",
		X"00",X"00",X"10",X"11",X"00",X"00",X"11",X"11",X"00",X"00",X"10",X"11",X"00",X"00",X"10",X"11",
		X"00",X"00",X"11",X"10",X"00",X"04",X"41",X"19",X"00",X"40",X"11",X"10",X"00",X"04",X"11",X"10",
		X"00",X"40",X"14",X"40",X"00",X"99",X"14",X"40",X"00",X"90",X"04",X"40",X"00",X"00",X"49",X"40",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"94",X"00",X"00",X"00",X"94",X"09",X"00",
		X"00",X"94",X"99",X"00",X"04",X"19",X"04",X"00",X"14",X"19",X"40",X"00",X"19",X"91",X"44",X"00",
		X"99",X"91",X"44",X"90",X"91",X"00",X"11",X"44",X"11",X"11",X"44",X"40",X"55",X"11",X"40",X"00",
		X"15",X"06",X"44",X"00",X"65",X"06",X"61",X"00",X"56",X"60",X"41",X"00",X"60",X"66",X"11",X"00",
		X"60",X"66",X"11",X"00",X"F0",X"66",X"01",X"00",X"66",X"00",X"66",X"99",X"00",X"66",X"11",X"14",
		X"FF",X"00",X"11",X"44",X"FF",X"00",X"00",X"44",X"00",X"0F",X"66",X"00",X"90",X"00",X"00",X"00",
		X"66",X"F0",X"11",X"00",X"06",X"00",X"09",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"01",X"11",X"00",X"00",X"00",X"91",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"33",X"00",X"00",X"33",X"30",X"00",X"00",X"36",X"39",X"00",X"00",X"36",X"36",X"00",
		X"00",X"36",X"39",X"00",X"00",X"93",X"90",X"90",X"00",X"33",X"39",X"00",X"00",X"61",X"39",X"00",
		X"00",X"36",X"46",X"00",X"00",X"11",X"66",X"00",X"00",X"66",X"61",X"00",X"00",X"66",X"41",X"00",
		X"00",X"44",X"63",X"00",X"00",X"33",X"16",X"00",X"00",X"36",X"13",X"00",X"00",X"36",X"11",X"00",
		X"00",X"99",X"31",X"90",X"00",X"39",X"33",X"30",X"00",X"39",X"13",X"39",X"00",X"90",X"13",X"03",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"99",X"00",X"90",X"00",X"93",X"00",X"00",
		X"00",X"96",X"90",X"00",X"00",X"96",X"99",X"00",X"01",X"66",X"99",X"00",X"06",X"36",X"61",X"00",
		X"00",X"66",X"61",X"09",X"99",X"66",X"11",X"99",X"96",X"66",X"19",X"39",X"66",X"66",X"19",X"69",
		X"66",X"61",X"16",X"99",X"00",X"6F",X"61",X"99",X"00",X"66",X"66",X"99",X"10",X"6F",X"11",X"90",
		X"69",X"FF",X"F3",X"90",X"90",X"FF",X"66",X"99",X"00",X"6F",X"66",X"99",X"00",X"4F",X"61",X"90",
		X"00",X"6F",X"66",X"90",X"00",X"FF",X"61",X"00",X"03",X"F6",X"66",X"90",X"06",X"66",X"16",X"99",
		X"66",X"61",X"96",X"99",X"99",X"11",X"11",X"99",X"99",X"31",X"99",X"99",X"90",X"93",X"99",X"99",
		X"00",X"39",X"99",X"90",X"00",X"90",X"19",X"99",X"00",X"00",X"19",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"90",X"90",X"00",X"09",X"90",X"99",X"00",X"99",X"99",X"09",X"00",X"39",X"00",X"00",
		X"00",X"39",X"09",X"99",X"00",X"36",X"99",X"90",X"00",X"36",X"99",X"00",X"01",X"61",X"93",X"09",
		X"03",X"39",X"99",X"33",X"00",X"69",X"11",X"99",X"09",X"31",X"99",X"33",X"03",X"63",X"99",X"96",
		X"00",X"16",X"61",X"39",X"00",X"63",X"13",X"99",X"00",X"06",X"99",X"39",X"00",X"03",X"13",X"93",
		X"00",X"63",X"39",X"33",X"00",X"66",X"99",X"93",X"00",X"34",X"93",X"99",X"00",X"36",X"19",X"09",
		X"03",X"36",X"11",X"00",X"00",X"33",X"11",X"30",X"30",X"33",X"99",X"30",X"00",X"33",X"69",X"33",
		X"61",X"13",X"99",X"99",X"30",X"39",X"19",X"99",X"30",X"19",X"99",X"39",X"00",X"39",X"99",X"99",
		X"00",X"91",X"93",X"63",X"00",X"09",X"99",X"90",X"00",X"00",X"30",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"90",X"00",X"00",
		X"00",X"90",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"93",X"00",X"00",X"19",X"99",X"00",
		X"00",X"19",X"33",X"00",X"00",X"11",X"33",X"09",X"00",X"39",X"33",X"93",X"00",X"99",X"99",X"33",
		X"00",X"16",X"93",X"33",X"00",X"11",X"33",X"93",X"09",X"99",X"93",X"99",X"39",X"61",X"99",X"00",
		X"90",X"93",X"93",X"00",X"93",X"63",X"69",X"00",X"39",X"19",X"39",X"33",X"99",X"11",X"33",X"93",
		X"03",X"91",X"93",X"90",X"93",X"61",X"03",X"00",X"93",X"69",X"93",X"00",X"93",X"96",X"93",X"99",
		X"39",X"99",X"39",X"33",X"09",X"01",X"39",X"33",X"09",X"99",X"13",X"39",X"03",X"09",X"99",X"99",
		X"00",X"09",X"96",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",
		X"00",X"30",X"99",X"00",X"00",X"33",X"39",X"00",X"00",X"33",X"33",X"00",X"00",X"33",X"39",X"33",
		X"00",X"33",X"93",X"00",X"00",X"33",X"39",X"90",X"00",X"33",X"93",X"33",X"00",X"33",X"99",X"33",
		X"00",X"33",X"93",X"33",X"00",X"33",X"93",X"30",X"00",X"93",X"33",X"00",X"00",X"99",X"93",X"00",
		X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"00",X"93",X"33",X"00",X"00",X"30",X"30",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"00",X"30",
		X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"03",
		X"00",X"50",X"00",X"30",X"00",X"03",X"05",X"90",X"00",X"35",X"33",X"00",X"00",X"03",X"33",X"00",
		X"00",X"F3",X"3F",X"30",X"00",X"F3",X"3F",X"90",X"00",X"F3",X"99",X"39",X"03",X"39",X"39",X"30",
		X"00",X"99",X"33",X"39",X"00",X"39",X"33",X"30",X"00",X"93",X"33",X"90",X"00",X"5F",X"35",X"00",
		X"00",X"5F",X"35",X"90",X"00",X"F0",X"35",X"33",X"00",X"39",X"95",X"00",X"00",X"3F",X"93",X"30",
		X"00",X"55",X"33",X"03",X"09",X"50",X"3F",X"00",X"53",X"53",X"3F",X"00",X"00",X"53",X"33",X"50",
		X"00",X"33",X"05",X"35",X"00",X"05",X"53",X"03",X"00",X"00",X"39",X"03",X"00",X"00",X"53",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"06",X"00",
		X"00",X"7F",X"04",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7F",X"01",X"00",
		X"00",X"7F",X"06",X"10",X"00",X"7F",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"06",X"00",
		X"00",X"FF",X"04",X"60",X"00",X"FF",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"F5",X"00",X"00",X"07",X"FF",X"01",X"00",
		X"07",X"FF",X"06",X"11",X"00",X"F5",X"00",X"06",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"07",X"F5",X"00",X"00",X"77",X"FF",X"00",X"00",X"77",X"FF",X"01",X"00",
		X"77",X"FF",X"06",X"11",X"07",X"F5",X"00",X"22",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"07",X"F5",X"00",X"00",X"77",X"FF",X"00",X"44",X"77",X"FF",X"06",X"00",
		X"77",X"FF",X"04",X"66",X"07",X"F5",X"00",X"22",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"40",X"00",
		X"00",X"04",X"64",X"00",X"00",X"00",X"60",X"00",X"00",X"44",X"94",X"00",X"00",X"00",X"64",X"00",
		X"00",X"00",X"04",X"00",X"00",X"04",X"44",X"00",X"00",X"90",X"04",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"40",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",X"0F",X"00",
		X"00",X"44",X"0F",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"F4",X"00",X"00",X"55",X"4F",X"00",
		X"00",X"44",X"64",X"00",X"00",X"44",X"64",X"00",X"00",X"44",X"64",X"00",X"00",X"F5",X"64",X"00",
		X"00",X"F0",X"64",X"00",X"00",X"F4",X"44",X"00",X"00",X"F5",X"44",X"00",X"00",X"3F",X"65",X"00",
		X"00",X"5F",X"60",X"00",X"00",X"00",X"40",X"00",X"00",X"05",X"46",X"00",X"00",X"00",X"40",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"5F",X"5F",X"00",
		X"00",X"44",X"5F",X"00",X"00",X"FF",X"FF",X"00",X"00",X"55",X"F4",X"00",X"00",X"55",X"4F",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"4F",X"64",X"00",X"00",X"FF",X"64",X"50",X"00",X"F5",X"6F",X"50",
		X"00",X"F5",X"44",X"50",X"00",X"F4",X"F4",X"00",X"00",X"F5",X"FF",X"00",X"00",X"3F",X"F5",X"00",
		X"00",X"5F",X"F5",X"00",X"00",X"F5",X"FF",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"0E",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"5F",X"55",X"00",
		X"03",X"5F",X"55",X"00",X"00",X"FF",X"53",X"00",X"00",X"55",X"35",X"00",X"00",X"55",X"3F",X"00",
		X"00",X"FF",X"5F",X"00",X"00",X"3F",X"FF",X"00",X"00",X"FF",X"FF",X"50",X"00",X"F5",X"FF",X"50",
		X"00",X"F5",X"F5",X"50",X"00",X"F5",X"F5",X"50",X"00",X"F5",X"FF",X"F0",X"00",X"3F",X"F5",X"00",
		X"00",X"5F",X"F5",X"50",X"00",X"55",X"FF",X"00",X"00",X"55",X"F5",X"00",X"00",X"55",X"FE",X"00",
		X"00",X"5F",X"E3",X"00",X"00",X"5F",X"05",X"00",X"00",X"F3",X"05",X"55",X"00",X"5F",X"00",X"55",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"55",X"EE",X"00",X"00",X"55",X"55",X"00",
		X"00",X"55",X"FF",X"00",X"00",X"F5",X"F5",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"55",X"00",
		X"00",X"5F",X"F5",X"00",X"00",X"EE",X"EF",X"00",X"0E",X"3F",X"3F",X"00",X"0E",X"FF",X"5F",X"00",
		X"0E",X"FF",X"5F",X"00",X"0E",X"5F",X"FF",X"00",X"0E",X"5F",X"55",X"00",X"0E",X"55",X"55",X"00",
		X"0E",X"35",X"F5",X"00",X"0E",X"F5",X"F5",X"00",X"00",X"35",X"55",X"00",X"00",X"F3",X"35",X"00",
		X"03",X"55",X"55",X"00",X"00",X"F5",X"55",X"35",X"03",X"35",X"55",X"33",X"00",X"53",X"FF",X"30",
		X"00",X"55",X"5F",X"00",X"00",X"F5",X"33",X"33",X"03",X"F5",X"EE",X"35",X"03",X"FF",X"00",X"F5",
		X"00",X"53",X"00",X"55",X"00",X"EE",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",X"04",X"00",
		X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"00",X"00",X"01",X"66",X"00",X"00",X"66",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"44",X"00",X"00",
		X"00",X"66",X"06",X"00",X"00",X"61",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"66",X"60",X"00",
		X"00",X"44",X"00",X"46",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"66",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"60",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"40",X"00",
		X"00",X"40",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"66",X"60",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"44",X"00",X"46",
		X"00",X"66",X"60",X"00",X"00",X"10",X"00",X"00",X"00",X"61",X"01",X"00",X"00",X"66",X"06",X"00",
		X"00",X"40",X"00",X"00",X"00",X"66",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"06",X"00",X"66",X"44",X"00",X"00",X"01",X"66",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"66",X"66",X"00",X"00",X"11",X"00",X"00",X"06",X"44",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"64",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"66",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"17",X"00",X"00",X"9F",X"77",X"00",X"00",
		X"09",X"07",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"90",X"90",X"00",X"11",X"09",X"00",
		X"00",X"11",X"99",X"00",X"00",X"F5",X"99",X"00",X"00",X"51",X"99",X"90",X"00",X"11",X"99",X"00",
		X"00",X"22",X"DD",X"99",X"00",X"7D",X"DD",X"90",X"00",X"77",X"DD",X"99",X"00",X"67",X"DA",X"90",
		X"00",X"77",X"DA",X"00",X"00",X"7D",X"DA",X"90",X"00",X"00",X"DA",X"09",X"00",X"00",X"AE",X"90",
		X"00",X"00",X"EE",X"09",X"00",X"00",X"EE",X"90",X"00",X"00",X"A0",X"90",X"00",X"00",X"DA",X"99",
		X"00",X"00",X"DA",X"9F",X"00",X"00",X"DD",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"0D",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"0D",X"99",X"00",X"00",X"0D",X"59",X"00",X"00",X"0D",X"55",
		X"00",X"00",X"DD",X"55",X"00",X"00",X"DD",X"94",X"00",X"00",X"AD",X"99",X"00",X"77",X"AA",X"90",
		X"00",X"77",X"7A",X"99",X"00",X"70",X"77",X"22",X"00",X"70",X"77",X"D2",X"00",X"00",X"D7",X"D2",
		X"00",X"00",X"D7",X"00",X"00",X"00",X"79",X"00",X"00",X"99",X"79",X"00",X"00",X"91",X"99",X"00",
		X"00",X"91",X"90",X"00",X"00",X"91",X"09",X"00",X"00",X"99",X"90",X"00",X"00",X"E9",X"09",X"00",
		X"00",X"E9",X"90",X"00",X"00",X"E5",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"69",X"99",X"0F",X"00",X"99",X"99",X"00",X"00",X"00",X"09",X"00",X"F0",X"0F",X"EE",
		X"0B",X"00",X"F9",X"EE",X"0B",X"AA",X"66",X"EE",X"0B",X"EB",X"A4",X"EE",X"0B",X"B5",X"64",X"00",
		X"00",X"05",X"49",X"EE",X"4B",X"05",X"9F",X"1E",X"04",X"01",X"FF",X"BB",X"0B",X"11",X"F0",X"00",
		X"BB",X"1F",X"FF",X"11",X"B0",X"1F",X"FF",X"F0",X"B0",X"1F",X"FF",X"55",X"A0",X"FF",X"1F",X"F5",
		X"A4",X"1F",X"FF",X"55",X"A6",X"1F",X"F1",X"55",X"B0",X"F1",X"FF",X"EB",X"0B",X"FF",X"10",X"EE",
		X"0F",X"66",X"BB",X"BE",X"F4",X"66",X"A9",X"EE",X"44",X"69",X"00",X"BE",X"40",X"00",X"90",X"EF",
		X"B0",X"00",X"60",X"FE",X"B0",X"AA",X"60",X"EF",X"BB",X"00",X"66",X"90",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"69",X"00",X"00",X"99",X"99",X"00",X"00",X"19",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"A0",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"F0",X"11",X"00",X"00",X"66",X"11",
		X"00",X"00",X"06",X"11",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"16",X"00",X"06",X"00",X"16",
		X"00",X"00",X"04",X"11",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"55",X"00",X"00",X"40",X"11",
		X"00",X"01",X"04",X"1F",X"00",X"00",X"66",X"FF",X"00",X"00",X"66",X"FF",X"00",X"00",X"14",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"B0",X"00",X"0F",X"66",X"3E",X"00",
		X"11",X"E6",X"0B",X"00",X"16",X"E0",X"03",X"00",X"61",X"00",X"00",X"00",X"46",X"06",X"11",X"00",
		X"66",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"F6",X"61",X"00",X"00",
		X"66",X"60",X"00",X"00",X"F5",X"11",X"0B",X"00",X"FF",X"BB",X"BB",X"00",X"FF",X"66",X"11",X"00",
		X"00",X"00",X"60",X"FF",X"00",X"00",X"44",X"FF",X"00",X"00",X"60",X"FF",X"00",X"00",X"00",X"1F",
		X"00",X"11",X"11",X"F1",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"66",X"00",X"00",X"66",X"16",
		X"00",X"00",X"60",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F6",X"44",X"EE",X"00",X"66",X"41",X"66",X"00",X"66",X"61",X"00",X"00",X"66",X"11",X"00",X"00",
		X"61",X"11",X"11",X"10",X"66",X"40",X"00",X"00",X"66",X"44",X"00",X"00",X"11",X"11",X"00",X"00",
		X"00",X"66",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"11",X"06",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"19",X"00",X"00",X"00",
		X"19",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"06",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"01",X"11",
		X"00",X"10",X"00",X"10",X"00",X"00",X"06",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"60",X"11",
		X"00",X"00",X"66",X"16",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"69",X"00",X"11",X"11",X"F1",
		X"00",X"00",X"00",X"1F",X"00",X"00",X"60",X"FF",X"00",X"00",X"44",X"FF",X"00",X"00",X"60",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"10",X"00",X"00",
		X"19",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"06",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"00",X"11",X"06",X"00",X"01",X"00",X"00",X"00",X"00",X"66",X"00",X"00",
		X"11",X"11",X"00",X"00",X"61",X"44",X"00",X"00",X"61",X"40",X"00",X"00",X"11",X"11",X"11",X"10",
		X"66",X"11",X"00",X"00",X"66",X"61",X"00",X"00",X"66",X"41",X"66",X"00",X"F6",X"44",X"EE",X"00",
		X"00",X"00",X"14",X"FF",X"00",X"00",X"66",X"FF",X"00",X"00",X"66",X"FF",X"00",X"01",X"04",X"1F",
		X"00",X"00",X"40",X"11",X"60",X"00",X"00",X"55",X"00",X"00",X"00",X"51",X"00",X"00",X"04",X"11",
		X"00",X"06",X"00",X"16",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"61",X"00",X"00",X"06",X"11",
		X"00",X"00",X"66",X"11",X"00",X"00",X"F0",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"66",X"11",X"00",X"FF",X"BB",X"0B",X"00",X"F5",X"11",X"00",X"00",X"66",X"60",X"00",X"00",
		X"F6",X"61",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"66",X"66",X"00",
		X"46",X"06",X"11",X"00",X"61",X"11",X"00",X"00",X"16",X"E0",X"03",X"00",X"11",X"E6",X"0B",X"00",
		X"0F",X"66",X"3E",X"00",X"99",X"00",X"B0",X"00",X"99",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",
		X"11",X"00",X"00",X"0A",X"66",X"11",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"16",X"00",X"00",
		X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"10",
		X"00",X"00",X"06",X"10",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"16",
		X"00",X"00",X"04",X"33",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"66",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"14",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"11",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A3",X"06",X"00",X"00",
		X"11",X"06",X"00",X"00",X"16",X"00",X"00",X"00",X"60",X"11",X"00",X"00",X"30",X"36",X"00",X"00",
		X"33",X"36",X"60",X"00",X"00",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"61",X"00",X"00",
		X"00",X"00",X"00",X"00",X"33",X"01",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"06",X"10",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"1F",
		X"00",X"00",X"11",X"30",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"36",X"00",X"00",X"66",X"33",
		X"00",X"00",X"60",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"10",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"33",X"66",X"00",X"00",X"61",X"33",X"00",X"00",X"11",X"00",X"00",
		X"00",X"11",X"01",X"00",X"00",X"40",X"00",X"00",X"33",X"44",X"00",X"00",X"03",X"11",X"00",X"00",
		X"03",X"63",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"33",X"00",X"00",X"00",X"00",X"00",
		X"63",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"03",X"00",X"10",X"00",X"19",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"AB",X"00",
		X"00",X"BB",X"00",X"A0",X"00",X"A0",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"42",X"99",X"11",
		X"00",X"77",X"99",X"FF",X"0B",X"55",X"FF",X"99",X"BA",X"55",X"FF",X"FF",X"BA",X"35",X"FF",X"99",
		X"AA",X"35",X"FF",X"9F",X"A5",X"55",X"FF",X"9F",X"A5",X"55",X"FF",X"9F",X"A5",X"55",X"FF",X"9F",
		X"A5",X"55",X"FF",X"9F",X"05",X"55",X"FF",X"9F",X"05",X"55",X"FF",X"9F",X"00",X"35",X"FF",X"9F",
		X"00",X"35",X"FF",X"99",X"B0",X"55",X"FF",X"FF",X"B0",X"55",X"FF",X"99",X"AB",X"77",X"99",X"FF",
		X"0B",X"42",X"99",X"11",X"0A",X"00",X"EE",X"BA",X"00",X"AA",X"AA",X"AA",X"00",X"0A",X"B0",X"00",
		X"00",X"00",X"A0",X"B0",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"AA",X"00",X"00",X"0A",
		X"00",X"AA",X"0A",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"55",X"FF",X"00",X"00",X"55",X"FF",X"F0",X"00",X"35",X"FF",X"99",
		X"00",X"35",X"FF",X"9F",X"00",X"55",X"FF",X"9F",X"0A",X"55",X"FF",X"9F",X"00",X"55",X"FF",X"9F",
		X"00",X"55",X"FF",X"9F",X"00",X"55",X"FF",X"9F",X"0A",X"55",X"FF",X"9F",X"0B",X"35",X"FF",X"9F",
		X"00",X"35",X"FF",X"99",X"00",X"55",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"0B",X"B0",X"00",X"0A",X"00",X"00",X"00",X"50",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"0B",X"00",X"BB",X"00",X"B0",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"A0",
		X"00",X"30",X"FF",X"00",X"0A",X"55",X"FF",X"00",X"0A",X"55",X"FF",X"00",X"00",X"55",X"FF",X"00",
		X"00",X"05",X"FF",X"00",X"00",X"00",X"FF",X"00",X"0A",X"00",X"FF",X"00",X"00",X"00",X"FF",X"B0",
		X"00",X"00",X"FF",X"B0",X"00",X"00",X"FF",X"BA",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"BB",X"00",X"0A",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",
		X"00",X"BB",X"00",X"00",X"00",X"0B",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"0A",X"00",X"B0",X"00",X"A0",X"00",X"B0",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"B0",X"0F",X"00",X"00",X"B0",X"00",X"A0",X"00",X"0B",X"00",X"A0",X"00",X"0B",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",
		X"00",X"00",X"F3",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"F3",X"00",X"00",X"01",X"93",X"00",
		X"00",X"01",X"93",X"00",X"00",X"01",X"F3",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",
		X"00",X"00",X"F3",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"F3",X"00",
		X"00",X"00",X"93",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"F3",X"00",
		X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"B0",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"0B",X"0B",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"0B",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",
		X"00",X"0B",X"00",X"00",X"B0",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"B0",X"00",X"0B",X"BB",X"B0",X"00",X"0B",X"BB",X"B0",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"B0",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"00",X"BB",
		X"BB",X"BB",X"0B",X"B0",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"0B",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"0B",X"0B",X"00",X"00",X"BB",X"BB",X"00",X"00",X"B0",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"0B",X"B0",
		X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"B0",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"00",X"B0",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"B0",X"00",X"0B",X"BB",X"B0",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"B0",X"00",
		X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"B0",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"99",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"92",X"22",X"22",X"92",X"99",X"99",X"99",X"92",X"92",X"22",X"22",X"92",
		X"22",X"97",X"22",X"22",X"22",X"97",X"22",X"22",X"22",X"77",X"22",X"22",X"22",X"79",X"22",X"22",
		X"22",X"7F",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",
		X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"22",
		X"22",X"FF",X"22",X"22",X"22",X"FF",X"22",X"92",X"22",X"99",X"2A",X"A9",X"22",X"FF",X"AA",X"AA",
		X"92",X"22",X"22",X"92",X"99",X"99",X"99",X"92",X"92",X"22",X"22",X"92",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"99",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"92",X"92",X"22",X"92",X"99",X"99",X"99",X"92",X"92",X"92",X"22",X"92",
		X"22",X"92",X"22",X"22",X"22",X"99",X"99",X"22",X"22",X"99",X"9E",X"22",X"22",X"E9",X"99",X"22",
		X"22",X"E9",X"99",X"22",X"22",X"99",X"99",X"22",X"22",X"99",X"99",X"22",X"22",X"E9",X"99",X"22",
		X"22",X"E9",X"99",X"22",X"22",X"E9",X"99",X"22",X"22",X"99",X"99",X"22",X"22",X"99",X"99",X"22",
		X"22",X"E9",X"99",X"22",X"22",X"EE",X"99",X"22",X"22",X"99",X"99",X"22",X"22",X"92",X"22",X"22",
		X"92",X"92",X"22",X"92",X"99",X"99",X"99",X"92",X"92",X"92",X"22",X"92",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"99",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"99",X"22",X"22",X"92",X"99",X"99",X"99",X"92",X"92",X"29",X"29",X"92",
		X"22",X"92",X"92",X"22",X"22",X"29",X"29",X"22",X"22",X"92",X"92",X"22",X"22",X"29",X"99",X"22",
		X"22",X"F5",X"99",X"22",X"22",X"F5",X"99",X"22",X"22",X"9F",X"55",X"22",X"22",X"9F",X"59",X"22",
		X"22",X"99",X"E9",X"22",X"22",X"5F",X"59",X"22",X"22",X"5F",X"E5",X"22",X"22",X"55",X"59",X"22",
		X"22",X"FF",X"92",X"22",X"22",X"F9",X"29",X"22",X"22",X"92",X"92",X"22",X"22",X"29",X"29",X"22",
		X"92",X"92",X"92",X"92",X"99",X"99",X"99",X"92",X"99",X"22",X"22",X"92",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",
		X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"90",
		X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",
		X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",
		X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"99",X"00",X"00",X"E5",X"55",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"09",X"FE",X"EE",X"00",X"9F",X"EE",X"99",X"00",X"FF",X"99",X"99",
		X"00",X"5F",X"EE",X"55",X"00",X"55",X"F5",X"99",X"00",X"F5",X"FF",X"EE",X"00",X"FF",X"FF",X"99",
		X"00",X"FF",X"EE",X"92",X"0F",X"FF",X"FF",X"92",X"FF",X"FF",X"FF",X"92",X"FF",X"EF",X"FF",X"92",
		X"FF",X"EF",X"FF",X"92",X"FF",X"FF",X"FF",X"92",X"0F",X"FF",X"FF",X"92",X"00",X"FF",X"FF",X"92",
		X"00",X"5F",X"FF",X"99",X"00",X"F5",X"FF",X"FF",X"00",X"FF",X"F5",X"99",X"00",X"FF",X"55",X"FF",
		X"00",X"FF",X"33",X"53",X"00",X"FF",X"55",X"33",X"00",X"5F",X"F5",X"55",X"00",X"00",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E5",X"99",X"99",X"00",X"55",X"55",X"55",X"00",
		X"FF",X"FF",X"FF",X"00",X"EE",X"FF",X"FF",X"00",X"EE",X"22",X"22",X"00",X"EF",X"44",X"42",X"00",
		X"F2",X"44",X"42",X"00",X"22",X"44",X"42",X"00",X"22",X"44",X"42",X"00",X"22",X"44",X"42",X"00",
		X"22",X"44",X"42",X"00",X"22",X"44",X"42",X"00",X"24",X"44",X"42",X"00",X"44",X"44",X"42",X"00",
		X"42",X"44",X"42",X"00",X"22",X"44",X"42",X"00",X"22",X"44",X"42",X"00",X"22",X"44",X"42",X"00",
		X"22",X"44",X"42",X"00",X"22",X"44",X"42",X"00",X"24",X"24",X"22",X"00",X"32",X"22",X"22",X"00",
		X"53",X"22",X"22",X"00",X"55",X"FF",X"FF",X"00",X"55",X"FF",X"FF",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"FF",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"EE",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"5E",
		X"00",X"99",X"99",X"3E",X"00",X"94",X"99",X"3E",X"00",X"49",X"95",X"3E",X"09",X"99",X"55",X"3E",
		X"09",X"99",X"55",X"3E",X"99",X"99",X"55",X"39",X"94",X"99",X"99",X"39",X"9A",X"AA",X"AA",X"39",
		X"94",X"AA",X"FF",X"39",X"9A",X"AA",X"FF",X"99",X"09",X"AA",X"FF",X"9E",X"09",X"AA",X"FF",X"9E",
		X"00",X"4A",X"AF",X"9E",X"00",X"A4",X"AA",X"9E",X"00",X"AA",X"AA",X"9E",X"00",X"9A",X"AA",X"FE",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"EE",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"E9",X"E9",X"00",X"00",X"E9",X"EE",X"00",X"00",X"E9",X"E5",X"00",X"00",
		X"E9",X"50",X"00",X"00",X"59",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",
		X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"99",X"99",X"C0",
		X"00",X"90",X"09",X"00",X"00",X"99",X"91",X"00",X"00",X"90",X"91",X"00",X"00",X"99",X"11",X"C0",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",
		X"00",X"99",X"11",X"00",X"00",X"90",X"91",X"00",X"00",X"99",X"91",X"00",X"00",X"90",X"09",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"FE",X"00",X"00",X"00",X"F3",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"F3",X"00",
		X"00",X"05",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"F3",X"50",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"F3",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"EF",X"50",X"00",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EF",X"00",
		X"00",X"00",X"99",X"05",X"00",X"00",X"EE",X"00",X"00",X"00",X"EF",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EF",X"F0",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"0C",X"99",X"C9",X"CC",X"C9",X"EB",X"0C",X"BB",X"65",X"CA",X"BE",X"9B",X"65",X"AA",X"AA",X"C9",
		X"65",X"BE",X"EB",X"BC",X"99",X"EB",X"BE",X"B9",X"5A",X"EB",X"BB",X"BB",X"5E",X"BB",X"BB",X"9B",
		X"5E",X"BB",X"BB",X"9A",X"FE",X"EE",X"B5",X"9A",X"F5",X"5F",X"BB",X"9A",X"FE",X"BB",X"5B",X"9A",
		X"5E",X"BB",X"B5",X"99",X"FE",X"BB",X"5B",X"9B",X"5E",X"BB",X"BF",X"BB",X"99",X"BB",X"FB",X"B9",
		X"65",X"96",X"BB",X"BC",X"65",X"BB",X"6F",X"CB",X"65",X"CC",X"BB",X"9B",X"CB",X"BB",X"0C",X"BB",
		X"0C",X"99",X"C9",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"99",X"00",X"77",X"99",X"99",X"00",X"77",X"DD",X"99",
		X"00",X"76",X"AD",X"99",X"00",X"07",X"DA",X"91",X"00",X"97",X"DD",X"19",X"04",X"19",X"AD",X"94",
		X"E6",X"11",X"7A",X"95",X"96",X"11",X"7A",X"55",X"E6",X"F1",X"7A",X"55",X"96",X"11",X"7A",X"95",
		X"04",X"17",X"7D",X"04",X"00",X"07",X"DD",X"10",X"00",X"97",X"DA",X"01",X"00",X"77",X"AD",X"00",
		X"00",X"76",X"D7",X"00",X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"99",X"99",X"39",X"0F",
		X"99",X"9A",X"E3",X"1F",X"99",X"99",X"99",X"91",X"F9",X"F9",X"99",X"10",X"99",X"99",X"99",X"41",
		X"0A",X"77",X"59",X"10",X"AA",X"AA",X"75",X"91",X"AA",X"AA",X"A7",X"10",X"AA",X"99",X"A5",X"90",
		X"AA",X"44",X"A7",X"90",X"AA",X"49",X"A7",X"90",X"AA",X"9A",X"AA",X"90",X"AA",X"94",X"AA",X"90",
		X"AA",X"49",X"AA",X"90",X"AA",X"94",X"AA",X"90",X"EA",X"9A",X"AE",X"90",X"AA",X"49",X"A5",X"90",
		X"EA",X"44",X"AE",X"90",X"AE",X"AE",X"E5",X"10",X"EE",X"EA",X"E5",X"91",X"EE",X"EE",X"59",X"10",
		X"99",X"99",X"99",X"41",X"F9",X"F9",X"99",X"10",X"99",X"99",X"99",X"91",X"99",X"9A",X"E3",X"1F",
		X"D9",X"D9",X"39",X"0F",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"03",X"10",X"00",X"00",X"99",X"01",X"00",X"00",
		X"EE",X"10",X"00",X"00",X"99",X"10",X"00",X"00",X"39",X"01",X"00",X"00",X"5E",X"10",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"5E",X"10",X"00",X"00",X"E9",X"01",X"00",X"00",X"33",X"10",X"00",X"00",
		X"99",X"10",X"00",X"00",X"99",X"01",X"00",X"00",X"33",X"10",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"07",X"60",X"00",X"00",X"11",X"01",X"00",X"00",X"70",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"70",X"60",X"00",X"00",X"11",X"01",X"00",X"00",X"07",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"09",X"90",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"99",X"99",X"99",X"00",X"AE",X"99",X"9E",X"00",X"5E",X"99",X"EE",X"00",X"E5",X"AE",X"99",
		X"00",X"5E",X"9A",X"9A",X"05",X"AA",X"A9",X"AF",X"05",X"99",X"9A",X"9A",X"05",X"97",X"99",X"99",
		X"05",X"9A",X"7A",X"7A",X"05",X"AA",X"5E",X"AE",X"05",X"AA",X"55",X"EA",X"05",X"AA",X"5E",X"AE",
		X"05",X"99",X"55",X"EA",X"05",X"99",X"5E",X"AE",X"05",X"E3",X"55",X"EE",X"05",X"EE",X"5E",X"EE",
		X"05",X"EE",X"55",X"EE",X"05",X"EE",X"5E",X"EE",X"05",X"EE",X"55",X"E5",X"05",X"9E",X"65",X"56",
		X"05",X"9E",X"AA",X"AA",X"05",X"99",X"DD",X"DD",X"05",X"EA",X"DD",X"DF",X"00",X"E5",X"DD",X"DD",
		X"00",X"5E",X"AA",X"AA",X"00",X"E5",X"EE",X"EA",X"00",X"EE",X"09",X"0E",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"AE",X"99",X"00",X"00",X"EA",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"9A",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"A9",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",
		X"AA",X"90",X"00",X"00",X"EA",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"11",X"FF",X"FF",X"09",X"11",X"55",X"55",X"09",X"11",X"9A",X"BB",X"09",X"11",X"9A",X"BB",
		X"02",X"11",X"9A",X"AB",X"00",X"19",X"99",X"AB",X"00",X"21",X"F9",X"AB",X"00",X"22",X"F9",X"AA",
		X"00",X"22",X"F9",X"99",X"00",X"22",X"F9",X"99",X"00",X"22",X"FF",X"FF",X"00",X"22",X"F9",X"AB",
		X"00",X"19",X"F9",X"9A",X"00",X"11",X"FF",X"9A",X"00",X"12",X"5F",X"9A",X"00",X"11",X"5F",X"9A",
		X"00",X"11",X"5F",X"9A",X"00",X"11",X"5F",X"99",X"00",X"11",X"5F",X"99",X"00",X"11",X"5F",X"FF",
		X"00",X"11",X"55",X"55",X"00",X"11",X"91",X"91",X"00",X"12",X"11",X"22",X"00",X"11",X"22",X"22",
		X"00",X"11",X"11",X"22",X"00",X"11",X"11",X"22",X"00",X"11",X"11",X"12",X"00",X"11",X"19",X"11",
		X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"0E",X"9E",X"EE",X"00",X"99",X"00",X"99",
		X"92",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",
		X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"29",X"99",X"39",X"22",
		X"92",X"22",X"92",X"29",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"33",X"22",X"32",X"32",X"99",X"99",X"39",X"33",
		X"33",X"33",X"33",X"33",X"33",X"33",X"13",X"33",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"91",X"12",X"22",X"22",X"22",X"11",X"12",X"11",
		X"21",X"91",X"11",X"11",X"91",X"11",X"11",X"11",X"91",X"11",X"11",X"11",X"21",X"11",X"11",X"11",
		X"91",X"11",X"19",X"19",X"91",X"11",X"92",X"29",X"21",X"11",X"99",X"99",X"22",X"22",X"99",X"99",
		X"00",X"99",X"33",X"99",X"00",X"3E",X"9E",X"EE",X"00",X"33",X"33",X"33",X"00",X"99",X"99",X"99",
		X"00",X"22",X"29",X"21",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"99",X"22",X"22",X"00",X"21",X"29",X"22",X"00",X"22",X"29",X"22",
		X"00",X"22",X"99",X"22",X"00",X"22",X"93",X"22",X"00",X"22",X"3E",X"22",X"00",X"99",X"3E",X"11",
		X"00",X"21",X"EE",X"99",X"00",X"22",X"FE",X"22",X"00",X"22",X"55",X"22",X"00",X"22",X"25",X"22",
		X"00",X"29",X"22",X"29",X"00",X"29",X"99",X"92",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"92",X"92",X"99",X"02",X"22",X"22",X"22",
		X"09",X"22",X"22",X"22",X"09",X"22",X"22",X"22",X"09",X"22",X"22",X"22",X"02",X"22",X"22",X"22",
		X"11",X"11",X"99",X"00",X"11",X"11",X"90",X"00",X"11",X"11",X"99",X"00",X"11",X"11",X"90",X"00",
		X"11",X"11",X"99",X"00",X"11",X"11",X"90",X"00",X"11",X"21",X"99",X"00",X"12",X"22",X"90",X"00",
		X"11",X"11",X"99",X"00",X"11",X"91",X"90",X"00",X"11",X"11",X"99",X"00",X"11",X"11",X"90",X"00",
		X"11",X"11",X"99",X"00",X"11",X"11",X"90",X"00",X"11",X"21",X"99",X"00",X"22",X"12",X"33",X"50",
		X"19",X"11",X"55",X"50",X"11",X"11",X"55",X"F0",X"11",X"11",X"55",X"F0",X"11",X"11",X"55",X"F0",
		X"11",X"11",X"35",X"F0",X"11",X"11",X"55",X"F0",X"22",X"22",X"35",X"F0",X"11",X"11",X"35",X"00",
		X"11",X"11",X"55",X"00",X"11",X"11",X"35",X"00",X"11",X"11",X"55",X"00",X"11",X"91",X"F9",X"00",
		X"99",X"99",X"90",X"00",X"EE",X"EE",X"90",X"00",X"EE",X"EE",X"90",X"00",X"E9",X"99",X"90",X"00",
		X"99",X"9F",X"90",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"90",X"00",X"22",X"22",X"99",X"00",
		X"22",X"22",X"90",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"90",X"00",X"99",X"9F",X"99",X"00",
		X"29",X"29",X"90",X"00",X"22",X"22",X"99",X"00",X"22",X"2F",X"90",X"00",X"22",X"2F",X"99",X"00",
		X"22",X"2F",X"90",X"00",X"22",X"2F",X"99",X"00",X"33",X"3F",X"90",X"00",X"99",X"FF",X"99",X"00",
		X"33",X"3F",X"90",X"00",X"33",X"3F",X"99",X"00",X"11",X"1F",X"90",X"00",X"11",X"1F",X"99",X"00",
		X"11",X"1F",X"90",X"00",X"11",X"19",X"99",X"00",X"11",X"19",X"90",X"00",X"12",X"29",X"99",X"00",
		X"11",X"12",X"90",X"00",X"11",X"11",X"99",X"00",X"11",X"11",X"90",X"00",X"11",X"11",X"99",X"00",
		X"11",X"11",X"90",X"00",X"12",X"11",X"99",X"00",X"22",X"11",X"90",X"00",X"11",X"22",X"99",X"00",
		X"19",X"99",X"90",X"00",X"EE",X"3E",X"90",X"00",X"33",X"33",X"90",X"00",X"99",X"99",X"90",X"00",
		X"11",X"91",X"F9",X"00",X"22",X"22",X"55",X"00",X"22",X"22",X"35",X"00",X"22",X"22",X"55",X"00",
		X"22",X"22",X"35",X"00",X"22",X"99",X"35",X"F0",X"21",X"12",X"55",X"F0",X"22",X"22",X"35",X"F0",
		X"22",X"22",X"55",X"F0",X"22",X"22",X"55",X"F0",X"22",X"22",X"55",X"F0",X"92",X"29",X"55",X"50",
		X"22",X"22",X"33",X"50",X"22",X"22",X"99",X"00",X"22",X"22",X"90",X"00",X"22",X"22",X"99",X"00",
		X"92",X"92",X"90",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"90",X"00",X"22",X"22",X"99",X"00",
		X"12",X"22",X"90",X"00",X"23",X"22",X"99",X"00",X"29",X"99",X"90",X"00",X"22",X"22",X"99",X"00",
		X"22",X"22",X"90",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"90",X"00",X"22",X"22",X"99",X"00",
		X"00",X"00",X"09",X"09",X"00",X"09",X"99",X"90",X"00",X"00",X"55",X"10",X"00",X"99",X"55",X"09",
		X"00",X"55",X"55",X"00",X"00",X"55",X"55",X"99",X"09",X"55",X"55",X"55",X"00",X"55",X"51",X"33",
		X"09",X"55",X"11",X"33",X"05",X"33",X"77",X"77",X"19",X"44",X"33",X"99",X"99",X"73",X"AB",X"33",
		X"55",X"33",X"BB",X"9D",X"0F",X"55",X"B9",X"9D",X"00",X"53",X"99",X"DD",X"00",X"33",X"99",X"DD",
		X"00",X"53",X"99",X"DD",X"00",X"F3",X"99",X"DD",X"03",X"FF",X"B9",X"9D",X"55",X"FF",X"BB",X"93",
		X"99",X"1F",X"AB",X"33",X"19",X"11",X"FF",X"FF",X"0F",X"55",X"11",X"11",X"00",X"55",X"11",X"55",
		X"00",X"55",X"51",X"55",X"00",X"55",X"55",X"FF",X"00",X"5F",X"55",X"00",X"00",X"FF",X"55",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"09",X"00",X"00",X"00",
		X"90",X"99",X"09",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"09",X"00",
		X"99",X"9F",X"00",X"00",X"FF",X"F5",X"90",X"00",X"59",X"55",X"09",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"99",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"99",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"09",X"00",X"F9",X"FF",X"90",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"55",X"FF",X"90",X"00",X"99",X"9F",X"00",X"00",X"F9",X"99",X"00",X"00",
		X"0F",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"91",X"00",X"09",X"99",X"16",X"00",
		X"90",X"96",X"66",X"00",X"09",X"61",X"10",X"60",X"99",X"69",X"10",X"00",X"99",X"99",X"09",X"00",
		X"99",X"9F",X"00",X"00",X"FF",X"F5",X"90",X"00",X"59",X"55",X"09",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"99",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"99",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"09",X"00",X"F9",X"FF",X"90",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"55",X"FF",X"90",X"00",X"99",X"9F",X"00",X"00",X"F9",X"99",X"00",X"00",
		X"0F",X"99",X"00",X"00",X"00",X"F9",X"60",X"60",X"00",X"0F",X"66",X"06",X"00",X"10",X"FF",X"00",
		X"00",X"61",X"11",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"09",X"00",X"00",X"00",
		X"90",X"99",X"09",X"00",X"09",X"96",X"60",X"00",X"99",X"99",X"66",X"00",X"99",X"99",X"69",X"00",
		X"99",X"9F",X"00",X"00",X"FF",X"F5",X"90",X"00",X"59",X"55",X"09",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"99",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"99",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"09",X"00",X"F9",X"FF",X"90",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"55",X"FF",X"90",X"00",X"99",X"9F",X"00",X"00",X"F9",X"99",X"00",X"00",
		X"0F",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"66",X"00",X"00",X"60",X"00",X"00",
		X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"17",X"00",X"00",X"00",X"77",X"00",X"00",X"00",
		X"71",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"F1",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"AE",X"99",X"00",X"00",X"EA",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"9A",X"99",X"00",X"00",X"A9",X"19",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"19",X"00",X"00",
		X"79",X"99",X"00",X"00",X"A9",X"19",X"00",X"00",X"79",X"99",X"00",X"00",X"A9",X"19",X"00",X"00",
		X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",X"79",X"99",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"79",X"19",X"00",X"00",X"A9",X"99",X"00",X"00",X"79",X"19",X"00",X"00",X"A9",X"99",X"00",X"00",
		X"A9",X"19",X"00",X"00",X"DD",X"99",X"00",X"00",X"DD",X"19",X"00",X"00",X"DD",X"99",X"00",X"00",
		X"AA",X"90",X"00",X"00",X"EA",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"11",X"11",
		X"00",X"00",X"17",X"11",X"00",X"09",X"72",X"21",X"00",X"21",X"29",X"29",X"00",X"11",X"92",X"92",
		X"00",X"77",X"99",X"99",X"00",X"22",X"44",X"49",X"00",X"22",X"44",X"42",X"00",X"22",X"49",X"49",
		X"00",X"22",X"22",X"42",X"0C",X"22",X"66",X"49",X"CC",X"22",X"29",X"42",X"CC",X"22",X"92",X"49",
		X"C6",X"22",X"29",X"42",X"EC",X"22",X"99",X"49",X"CC",X"22",X"99",X"42",X"6C",X"92",X"99",X"49",
		X"CC",X"29",X"99",X"42",X"66",X"92",X"F6",X"49",X"06",X"39",X"77",X"42",X"00",X"93",X"44",X"49",
		X"00",X"90",X"44",X"49",X"00",X"29",X"92",X"92",X"00",X"12",X"29",X"29",X"00",X"11",X"92",X"92",
		X"00",X"17",X"99",X"99",X"00",X"06",X"22",X"21",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"12",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"99",X"00",X"00",X"11",X"92",X"99",X"00",
		X"11",X"21",X"92",X"00",X"12",X"11",X"12",X"00",X"22",X"21",X"11",X"00",X"22",X"92",X"91",X"00",
		X"22",X"92",X"29",X"90",X"27",X"92",X"92",X"90",X"07",X"92",X"99",X"00",X"27",X"22",X"29",X"90",
		X"27",X"92",X"99",X"00",X"27",X"22",X"29",X"90",X"27",X"22",X"99",X"00",X"22",X"22",X"29",X"90",
		X"22",X"22",X"99",X"00",X"22",X"22",X"29",X"90",X"22",X"22",X"99",X"00",X"22",X"22",X"29",X"00",
		X"22",X"22",X"99",X"00",X"22",X"22",X"29",X"00",X"22",X"22",X"92",X"00",X"24",X"22",X"20",X"00",
		X"22",X"92",X"91",X"00",X"22",X"29",X"11",X"00",X"92",X"99",X"11",X"00",X"99",X"22",X"10",X"00",
		X"11",X"11",X"00",X"00",X"11",X"12",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",
		X"00",X"05",X"05",X"00",X"00",X"55",X"50",X"00",X"00",X"55",X"55",X"00",X"55",X"0F",X"00",X"00",
		X"55",X"55",X"55",X"00",X"55",X"50",X"55",X"00",X"00",X"50",X"55",X"00",X"00",X"05",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"50",X"00",X"00",X"50",X"05",X"00",X"FF",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"50",X"50",X"05",X"05",X"00",X"55",X"00",X"55",X"50",X"50",X"00",X"55",X"00",X"F5",
		X"00",X"50",X"50",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"50",X"00",X"00",X"F5",X"50",X"00",
		X"00",X"55",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"5F",X"50",X"00",X"00",X"F5",X"55",X"00",
		X"00",X"55",X"50",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"55",X"00",X"00",X"55",X"50",X"00",
		X"00",X"55",X"50",X"00",X"00",X"05",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"55",X"11",X"50",X"00",X"95",X"11",X"55",X"00",
		X"91",X"11",X"55",X"00",X"99",X"51",X"55",X"00",X"19",X"55",X"55",X"00",X"11",X"55",X"55",X"00",
		X"11",X"53",X"55",X"00",X"51",X"33",X"55",X"00",X"51",X"55",X"11",X"00",X"55",X"F5",X"11",X"50",
		X"55",X"F5",X"11",X"11",X"F5",X"5F",X"11",X"99",X"F5",X"F5",X"11",X"99",X"F5",X"F9",X"F1",X"99",
		X"F5",X"F9",X"BF",X"99",X"FF",X"F9",X"BB",X"09",X"0F",X"F9",X"9B",X"09",X"0F",X"F9",X"99",X"00",
		X"0F",X"FF",X"19",X"F0",X"00",X"1F",X"11",X"50",X"00",X"11",X"59",X"5F",X"00",X"11",X"99",X"5F",
		X"00",X"11",X"99",X"55",X"00",X"11",X"9D",X"25",X"00",X"11",X"9D",X"15",X"00",X"19",X"09",X"12",
		X"11",X"20",X"F9",X"99",X"11",X"11",X"FF",X"99",X"19",X"11",X"FF",X"FF",X"19",X"55",X"F9",X"0F",
		X"19",X"55",X"99",X"00",X"09",X"FF",X"9F",X"99",X"09",X"00",X"F9",X"99",X"00",X"90",X"39",X"FF",
		X"00",X"09",X"3F",X"1F",X"00",X"90",X"13",X"11",X"00",X"00",X"11",X"31",X"00",X"00",X"F1",X"31",
		X"00",X"00",X"F1",X"F3",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"F9",X"F9",
		X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"09",X"00",X"00",X"F9",X"90",X"00",X"00",X"F9",X"09",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"99",X"90",X"DD",X"00",X"09",X"00",X"BB",X"00",X"09",X"00",X"99",
		X"00",X"09",X"09",X"99",X"00",X"49",X"D9",X"99",X"00",X"B4",X"DD",X"99",X"00",X"BB",X"DD",X"99",
		X"00",X"FB",X"99",X"99",X"99",X"BF",X"99",X"99",X"9D",X"99",X"BB",X"99",X"29",X"94",X"BB",X"99",
		X"22",X"4F",X"BB",X"99",X"22",X"FF",X"FB",X"99",X"22",X"FF",X"BB",X"99",X"22",X"FF",X"FB",X"99",
		X"22",X"FF",X"BB",X"99",X"22",X"99",X"FB",X"99",X"22",X"49",X"BF",X"99",X"2A",X"F4",X"FB",X"99",
		X"AB",X"FF",X"BF",X"99",X"9B",X"FF",X"F9",X"99",X"0A",X"FF",X"9A",X"99",X"00",X"F9",X"9A",X"99",
		X"00",X"94",X"AA",X"99",X"00",X"4B",X"99",X"99",X"00",X"99",X"09",X"99",X"00",X"09",X"00",X"99",
		X"00",X"09",X"00",X"DD",X"00",X"99",X"90",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"D9",X"A9",X"00",X"AA",
		X"9B",X"DB",X"9A",X"A9",X"BD",X"BD",X"BD",X"99",X"BB",X"BB",X"BB",X"BB",X"5F",X"FF",X"FF",X"BF",
		X"B5",X"55",X"B5",X"BB",X"BB",X"BB",X"BB",X"AA",X"DB",X"DB",X"AA",X"BB",X"DD",X"AA",X"00",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"DD",X"90",X"00",X"00",X"9D",X"90",X"00",X"00",X"B9",X"99",X"00",
		X"00",X"BB",X"99",X"00",X"00",X"BB",X"99",X"D0",X"00",X"BB",X"99",X"DD",X"00",X"BB",X"49",X"BD",
		X"00",X"BB",X"49",X"0D",X"00",X"FB",X"4B",X"0B",X"00",X"B4",X"4B",X"00",X"00",X"F4",X"BB",X"00",
		X"00",X"44",X"BB",X"0E",X"00",X"F4",X"BB",X"90",X"00",X"FF",X"BB",X"99",X"00",X"FF",X"BB",X"99",
		X"00",X"FF",X"FB",X"99",X"00",X"44",X"BB",X"9A",X"00",X"BB",X"FB",X"9B",X"09",X"BB",X"BB",X"9B",
		X"00",X"99",X"FB",X"BB",X"00",X"00",X"A9",X"F9",X"00",X"00",X"AA",X"BF",X"00",X"00",X"A9",X"9F",
		X"00",X"99",X"99",X"B9",X"00",X"09",X"00",X"BB",X"00",X"00",X"99",X"EB",X"00",X"00",X"99",X"0E",
		X"00",X"00",X"B9",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0F",X"00",
		X"D0",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"D0",X"00",X"00",
		X"BF",X"DD",X"00",X"00",X"BB",X"BD",X"00",X"00",X"DB",X"BB",X"00",X"00",X"0D",X"FB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BB",X"00",X"D0",X"00",X"DB",X"D0",X"DD",
		X"00",X"DD",X"BD",X"BD",X"00",X"00",X"BB",X"BD",X"00",X"00",X"FB",X"A0",X"00",X"00",X"BF",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"F0",X"00",X"00",X"0B",X"00",X"00",X"00",X"AB",X"00",
		X"00",X"00",X"AB",X"00",X"00",X"00",X"AA",X"BB",X"00",X"00",X"0A",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"D9",X"90",X"00",
		X"22",X"DD",X"90",X"00",X"22",X"FB",X"09",X"00",X"22",X"FF",X"09",X"00",X"2F",X"FF",X"09",X"00",
		X"FB",X"9F",X"00",X"00",X"AF",X"F9",X"00",X"00",X"AA",X"9F",X"00",X"00",X"44",X"49",X"00",X"00",
		X"FF",X"F4",X"00",X"00",X"FF",X"F9",X"90",X"00",X"9F",X"94",X"90",X"00",X"9F",X"44",X"90",X"00",
		X"99",X"4F",X"99",X"00",X"44",X"FB",X"90",X"00",X"B4",X"BB",X"90",X"00",X"BB",X"FB",X"90",X"00",
		X"BB",X"BB",X"90",X"00",X"BB",X"BB",X"90",X"90",X"9B",X"BB",X"90",X"D0",X"9A",X"BB",X"90",X"D9",
		X"09",X"BB",X"00",X"D9",X"00",X"AB",X"09",X"D9",X"00",X"BA",X"99",X"BD",X"00",X"9B",X"B9",X"B0",
		X"00",X"9B",X"B9",X"00",X"90",X"B9",X"BB",X"00",X"90",X"EB",X"B9",X"00",X"99",X"00",X"9A",X"00",
		X"09",X"09",X"AA",X"00",X"00",X"99",X"BB",X"00",X"00",X"99",X"0B",X"00",X"00",X"99",X"FB",X"00",
		X"00",X"99",X"BF",X"00",X"00",X"99",X"BF",X"00",X"00",X"90",X"BB",X"00",X"00",X"00",X"DB",X"00",
		X"00",X"00",X"DB",X"00",X"00",X"00",X"AD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BD",
		X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"AB",X"00",X"00",X"0A",X"DB",X"00",X"00",X"AA",X"DD",
		X"00",X"00",X"0A",X"9D",X"00",X"00",X"09",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0B",X"00",X"BB",X"0B",X"00",X"00",X"99",X"0B",X"00",X"00",X"D9",X"0B",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"BD",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"BD",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"D9",X"00",
		X"00",X"00",X"BD",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"D0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"FB",X"AA",X"D0",X"00",X"BB",X"AA",X"D0",X"00",X"BB",X"AA",X"D0",
		X"00",X"AB",X"AA",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"00",
		X"00",X"90",X"22",X"00",X"00",X"00",X"2A",X"00",X"00",X"0A",X"2A",X"00",X"00",X"AA",X"AD",X"00",
		X"00",X"AB",X"99",X"00",X"00",X"AB",X"B9",X"00",X"00",X"BB",X"B9",X"09",X"00",X"AA",X"BB",X"09",
		X"00",X"44",X"4B",X"99",X"00",X"FF",X"44",X"09",X"00",X"FF",X"49",X"09",X"00",X"9F",X"F4",X"09",
		X"00",X"49",X"F4",X"09",X"00",X"94",X"F4",X"09",X"00",X"A9",X"99",X"09",X"00",X"A9",X"44",X"09",
		X"00",X"A9",X"FB",X"09",X"00",X"A9",X"BF",X"99",X"00",X"A9",X"FB",X"00",X"00",X"AA",X"BB",X"00",
		X"00",X"AA",X"BB",X"00",X"05",X"AA",X"BB",X"00",X"09",X"9A",X"BA",X"00",X"09",X"9A",X"BB",X"00",
		X"0B",X"99",X"BA",X"0B",X"09",X"09",X"BB",X"0B",X"0B",X"00",X"99",X"0B",X"09",X"99",X"99",X"9B",
		X"0B",X"99",X"BB",X"9B",X"09",X"99",X"59",X"9B",X"0B",X"99",X"B9",X"9B",X"09",X"99",X"59",X"9B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"BD",
		X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"40",X"00",X"00",X"66",X"00",X"00",X"46",X"66",X"00",
		X"00",X"60",X"66",X"00",X"00",X"40",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"06",X"00",X"00",X"66",X"00",X"00",X"46",X"44",X"00",X"00",X"60",X"44",X"00",
		X"00",X"60",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"04",X"66",X"00",X"00",X"06",X"66",X"60",
		X"00",X"00",X"44",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"04",X"66",X"00",X"00",X"66",X"66",X"40",X"00",X"06",X"64",X"04",X"00",X"00",X"66",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"46",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"60",X"00",X"46",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"60",X"00",
		X"00",X"00",X"00",X"04",X"64",X"00",X"66",X"00",X"06",X"46",X"44",X"00",X"06",X"60",X"44",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"06",X"66",X"40",
		X"00",X"00",X"44",X"00",X"00",X"04",X"04",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"64",X"66",X"00",X"00",X"66",X"66",X"60",X"00",X"06",X"64",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"46",X"00",
		X"00",X"40",X"66",X"00",X"00",X"64",X"66",X"44",X"04",X"66",X"66",X"40",X"06",X"66",X"66",X"00",
		X"66",X"60",X"66",X"00",X"00",X"00",X"66",X"00",X"40",X"06",X"06",X"00",X"64",X"66",X"66",X"00",
		X"66",X"00",X"06",X"04",X"66",X"00",X"66",X"00",X"06",X"46",X"44",X"00",X"00",X"66",X"64",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"06",X"66",X"00",X"40",X"00",X"44",X"40",
		X"64",X"00",X"66",X"60",X"66",X"64",X"66",X"00",X"06",X"66",X"66",X"00",X"00",X"66",X"66",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"40",X"06",X"06",X"64",X"00",X"00",X"00",X"66",X"00",
		X"00",X"04",X"40",X"00",X"00",X"66",X"60",X"00",X"00",X"46",X"06",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"40",X"40",X"66",X"06",X"66",X"04",X"06",X"66",X"64",X"00",X"66",X"40",X"06",X"00",X"66",X"00",
		X"66",X"00",X"66",X"00",X"00",X"06",X"60",X"00",X"40",X"00",X"06",X"00",X"64",X"00",X"66",X"40",
		X"66",X"00",X"06",X"66",X"66",X"00",X"66",X"66",X"06",X"40",X"44",X"00",X"00",X"40",X"64",X"00",
		X"00",X"60",X"66",X"00",X"06",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"40",X"00",X"44",X"40",
		X"64",X"00",X"66",X"60",X"66",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"06",X"06",X"00",X"46",X"00",X"00",X"66",X"66",X"00",X"64",X"00",X"00",X"00",X"66",X"00",
		X"00",X"04",X"40",X"00",X"00",X"66",X"60",X"40",X"00",X"40",X"06",X"60",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"0A",X"0F",X"00",X"A0",X"A0",X"F0",X"00",X"0A",X"FA",X"00",X"A0",X"A0",X"0F",X"0F",
		X"0A",X"F0",X"00",X"00",X"A0",X"00",X"00",X"00",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"A0",X"A0",X"00",X"0A",X"00",X"00",X"00",X"A0",X"A0",X"00",X"00",X"FF",X"0A",X"00",X"00",
		X"00",X"A0",X"0A",X"00",X"0F",X"00",X"A0",X"00",X"F0",X"FA",X"0A",X"A0",X"00",X"0F",X"00",X"00",
		X"00",X"F0",X"F0",X"0A",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"A0",X"0A",X"A0",X"00",X"0A",X"A0",X"0F",
		X"00",X"A0",X"0A",X"F0",X"A0",X"0A",X"00",X"00",X"0A",X"F0",X"00",X"00",X"F0",X"0F",X"F0",X"00",
		X"A0",X"A0",X"A0",X"00",X"0A",X"00",X"00",X"00",X"F0",X"A0",X"00",X"00",X"0F",X"0A",X"A0",X"00",
		X"00",X"F0",X"0A",X"A0",X"00",X"0F",X"A0",X"00",X"00",X"00",X"0F",X"A0",X"00",X"0F",X"F0",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"F0",X"0F",
		X"00",X"00",X"0F",X"00",X"00",X"F0",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"F0",X"FF",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"F0",X"0F",X"FF",X"00",X"F0",X"00",X"0F",X"0F",X"00",X"00",X"F0",X"0F",
		X"00",X"00",X"FF",X"00",X"00",X"F0",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"0F",X"FF",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"0F",X"0F",X"FF",X"00",X"00",X"F0",X"FF",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"0F",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"FF",X"00",X"F0",X"00",X"0F",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"F0",X"0F",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"F0",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"39",X"30",X"90",X"00",X"B3",X"B3",X"30",X"00",X"BB",X"BB",X"B0",
		X"00",X"5F",X"55",X"50",X"00",X"B3",X"B3",X"30",X"00",X"39",X"30",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"39",X"30",X"90",X"00",X"B3",X"B3",X"30",X"00",X"B5",X"55",X"50",
		X"00",X"5F",X"55",X"50",X"00",X"B3",X"B3",X"30",X"00",X"39",X"30",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"50",X"00",X"00",
		X"00",X"05",X"00",X"00",X"50",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"93",X"00",X"00",X"30",X"30",X"09",X"00",X"00",X"00",X"90",X"0F",
		X"05",X"05",X"35",X"50",X"30",X"30",X"03",X"00",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"93",X"00",X"00",X"30",X"30",X"09",X"00",X"00",X"00",X"90",X"50",
		X"05",X"05",X"35",X"00",X"30",X"30",X"03",X"F0",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"E9",X"99",X"00",X"00",X"D9",X"99",X"00",X"09",X"99",X"99",
		X"00",X"9D",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"DD",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"DD",X"EE",X"55",X"00",X"99",X"B5",X"99",X"00",X"DD",X"5B",X"EE",X"09",X"99",X"B5",X"99",
		X"9D",X"DD",X"99",X"99",X"99",X"99",X"F5",X"9A",X"DD",X"D9",X"5F",X"99",X"99",X"9E",X"FF",X"9A",
		X"AA",X"9A",X"5F",X"99",X"AB",X"A5",X"FF",X"9A",X"BA",X"BA",X"5F",X"99",X"0B",X"AB",X"55",X"9A",
		X"0A",X"BA",X"5B",X"99",X"00",X"AB",X"B5",X"FF",X"00",X"BA",X"5B",X"99",X"00",X"AB",X"55",X"55",
		X"00",X"BA",X"99",X"99",X"00",X"AB",X"55",X"99",X"00",X"BA",X"BA",X"AA",X"00",X"AB",X"AB",X"BB",
		X"00",X"0B",X"BA",X"AA",X"00",X"00",X"AB",X"BB",X"00",X"00",X"BA",X"BA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"9D",X"9D",X"00",
		X"99",X"DD",X"DD",X"00",X"99",X"9D",X"D9",X"00",X"99",X"BB",X"BB",X"00",X"99",X"DD",X"DD",X"00",
		X"99",X"BB",X"BB",X"00",X"9E",X"DD",X"DD",X"00",X"EA",X"BB",X"BB",X"00",X"AE",X"DD",X"DD",X"00",
		X"EA",X"BB",X"BB",X"00",X"AE",X"BD",X"DB",X"00",X"AA",X"BB",X"BB",X"00",X"A9",X"BB",X"BB",X"00",
		X"9A",X"BB",X"AB",X"00",X"AA",X"BB",X"BB",X"00",X"9A",X"AB",X"AB",X"00",X"A9",X"BB",X"BB",X"00",
		X"99",X"AA",X"AA",X"00",X"99",X"BB",X"BB",X"00",X"99",X"AA",X"AA",X"00",X"59",X"BB",X"BB",X"00",
		X"55",X"AA",X"AA",X"00",X"55",X"BB",X"BB",X"00",X"AA",X"AA",X"AA",X"00",X"BB",X"BA",X"AA",X"00",
		X"AA",X"AA",X"AA",X"00",X"AB",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"9A",X"9A",X"00",X"AB",X"AB",X"AB",X"00",X"BD",X"BD",X"BD",X"00",X"BB",X"BB",X"BB",
		X"00",X"5B",X"5B",X"5B",X"00",X"BA",X"BA",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"BA",X"BA",X"BA",
		X"00",X"AB",X"AB",X"AB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"AB",X"AB",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"FF",X"00",X"FF",X"FF",X"00",X"00",X"F0",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"0F",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"0F",X"F0",X"00",X"00",X"0F",X"F5",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"0F",X"F0",X"00",
		X"00",X"0F",X"00",X"00",X"0F",X"00",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"FF",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"00",X"FF",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"F0",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"F0",X"F0",X"00",X"F0",X"00",X"00",X"00",
		X"0F",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"F0",X"0F",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"F0",X"00",X"00",X"99",X"FF",X"00",X"99",X"95",X"AA",
		X"00",X"99",X"55",X"03",X"00",X"99",X"55",X"93",X"00",X"95",X"55",X"95",X"00",X"99",X"33",X"93",
		X"00",X"95",X"77",X"77",X"00",X"11",X"33",X"99",X"00",X"44",X"33",X"BB",X"00",X"57",X"33",X"99",
		X"00",X"15",X"5A",X"99",X"00",X"95",X"5A",X"99",X"00",X"55",X"AA",X"99",X"00",X"FF",X"AA",X"99",
		X"00",X"9F",X"99",X"99",X"00",X"19",X"99",X"19",X"00",X"51",X"99",X"19",X"00",X"99",X"99",X"59",
		X"00",X"99",X"9F",X"FF",X"09",X"99",X"11",X"11",X"00",X"99",X"55",X"95",X"00",X"99",X"55",X"95",
		X"00",X"99",X"55",X"93",X"00",X"00",X"55",X"93",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"19",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",
		X"90",X"99",X"00",X"00",X"59",X"FF",X"03",X"00",X"55",X"00",X"30",X"00",X"35",X"33",X"03",X"00",
		X"39",X"33",X"30",X"00",X"99",X"33",X"33",X"00",X"11",X"33",X"30",X"F0",X"59",X"93",X"0F",X"F0",
		X"59",X"6F",X"0F",X"00",X"55",X"66",X"00",X"F0",X"55",X"9F",X"FF",X"F0",X"55",X"9F",X"0F",X"00",
		X"55",X"99",X"FF",X"00",X"59",X"FF",X"00",X"00",X"59",X"99",X"00",X"00",X"14",X"11",X"F0",X"00",
		X"F5",X"FF",X"0F",X"00",X"5F",X"F9",X"0F",X"00",X"5F",X"0F",X"00",X"00",X"F0",X"00",X"FF",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"0F",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"FF",X"F0",X"00",X"0F",X"F0",X"0F",X"00",X"F0",X"00",X"00",X"00",X"09",X"55",X"00",
		X"00",X"99",X"99",X"00",X"00",X"59",X"55",X"19",X"00",X"59",X"55",X"99",X"00",X"99",X"33",X"99",
		X"00",X"95",X"47",X"77",X"00",X"91",X"93",X"39",X"00",X"94",X"33",X"BB",X"00",X"59",X"33",X"99",
		X"00",X"19",X"55",X"99",X"00",X"19",X"55",X"99",X"00",X"95",X"5A",X"99",X"00",X"9F",X"5A",X"99",
		X"00",X"19",X"95",X"99",X"00",X"11",X"99",X"99",X"00",X"95",X"99",X"99",X"00",X"44",X"99",X"19",
		X"00",X"11",X"91",X"11",X"00",X"95",X"41",X"11",X"00",X"99",X"55",X"15",X"00",X"99",X"55",X"59",
		X"00",X"99",X"55",X"19",X"00",X"90",X"95",X"19",X"00",X"00",X"9F",X"19",X"00",X"00",X"9F",X"11",
		X"00",X"00",X"99",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"90",X"00",X"0F",
		X"00",X"90",X"F0",X"00",X"55",X"00",X"F0",X"0F",X"55",X"F0",X"03",X"F0",X"33",X"00",X"00",X"FF",
		X"33",X"50",X"33",X"00",X"39",X"00",X"30",X"FF",X"41",X"0F",X"30",X"0F",X"95",X"00",X"30",X"0F",
		X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"0F",X"55",X"00",X"0F",X"0F",X"55",X"F0",X"00",X"00",
		X"55",X"F0",X"0F",X"F0",X"F5",X"F0",X"00",X"00",X"95",X"99",X"00",X"F0",X"11",X"11",X"0F",X"00",
		X"FF",X"FF",X"00",X"FF",X"F5",X"FF",X"00",X"0F",X"55",X"00",X"00",X"00",X"5F",X"E0",X"F0",X"0F",
		X"F0",X"90",X"F0",X"0F",X"00",X"90",X"0F",X"00",X"0F",X"F0",X"F0",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"0F",X"0F",X"00",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"FF",X"F0",X"0F",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"99",
		X"0F",X"05",X"33",X"99",X"00",X"99",X"47",X"77",X"00",X"91",X"93",X"39",X"0F",X"44",X"33",X"BB",
		X"F0",X"55",X"33",X"00",X"F0",X"11",X"55",X"00",X"00",X"15",X"55",X"00",X"FF",X"55",X"5A",X"00",
		X"00",X"FF",X"5A",X"99",X"00",X"1F",X"99",X"99",X"00",X"91",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"49",X"99",X"99",X"00",X"11",X"99",X"FF",X"00",X"95",X"49",X"19",X"00",X"99",X"55",X"F9",
		X"00",X"99",X"55",X"F9",X"00",X"99",X"55",X"99",X"00",X"90",X"95",X"99",X"00",X"00",X"99",X"99",
		X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"91",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"55",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"50",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"F5",X"F0",X"00",X"00",X"95",X"0F",X"00",X"00",
		X"11",X"00",X"0F",X"00",X"FF",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"5F",X"00",X"F0",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"0F",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"0F",X"0F",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"F0",X"00",X"01",X"00",X"0F",X"00",X"00",X"F0",X"F0",X"55",X"00",X"FF",X"00",X"95",X"10",
		X"F0",X"99",X"53",X"11",X"00",X"00",X"34",X"77",X"00",X"90",X"43",X"99",X"F0",X"04",X"93",X"BB",
		X"0F",X"59",X"33",X"90",X"00",X"FF",X"33",X"00",X"0F",X"81",X"35",X"00",X"F0",X"11",X"55",X"00",
		X"00",X"91",X"55",X"00",X"00",X"99",X"39",X"00",X"00",X"93",X"39",X"00",X"0F",X"95",X"F9",X"00",
		X"00",X"94",X"FF",X"99",X"00",X"00",X"11",X"FF",X"00",X"00",X"04",X"51",X"00",X"00",X"00",X"5F",
		X"00",X"00",X"55",X"55",X"0F",X"00",X"99",X"55",X"0F",X"F9",X"00",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",
		X"0F",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"F0",X"00",X"30",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",
		X"95",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"F0",X"00",X"00",
		X"00",X"33",X"99",X"00",X"00",X"FF",X"90",X"00",X"09",X"55",X"39",X"00",X"99",X"55",X"F3",X"00",
		X"99",X"55",X"FF",X"00",X"99",X"11",X"FF",X"09",X"F5",X"11",X"55",X"09",X"FF",X"11",X"55",X"01",
		X"FF",X"FF",X"55",X"99",X"FF",X"99",X"91",X"99",X"9F",X"99",X"91",X"99",X"91",X"9F",X"99",X"99",
		X"99",X"5F",X"99",X"33",X"99",X"5F",X"BB",X"53",X"09",X"95",X"99",X"5F",X"50",X"9F",X"99",X"55",
		X"55",X"FF",X"99",X"55",X"F5",X"FF",X"99",X"15",X"9F",X"11",X"99",X"15",X"99",X"11",X"99",X"19",
		X"99",X"11",X"99",X"F1",X"09",X"51",X"B9",X"99",X"00",X"55",X"1F",X"99",X"00",X"55",X"11",X"99",
		X"00",X"5F",X"91",X"99",X"00",X"55",X"95",X"99",X"00",X"FF",X"95",X"99",X"00",X"FF",X"95",X"99",
		X"00",X"9F",X"95",X"F9",X"00",X"FF",X"99",X"F9",X"00",X"00",X"99",X"FF",X"00",X"00",X"90",X"FF",
		X"9F",X"10",X"00",X"00",X"99",X"10",X"00",X"00",X"99",X"F1",X"00",X"00",X"99",X"91",X"99",X"00",
		X"90",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"55",X"39",X"00",
		X"00",X"95",X"99",X"00",X"00",X"F9",X"F9",X"00",X"00",X"11",X"11",X"30",X"00",X"11",X"99",X"F0",
		X"00",X"99",X"FF",X"00",X"00",X"5F",X"99",X"00",X"00",X"F9",X"FF",X"00",X"00",X"59",X"FF",X"00",
		X"00",X"F9",X"99",X"00",X"00",X"F9",X"FF",X"00",X"00",X"99",X"99",X"F0",X"00",X"94",X"11",X"00",
		X"00",X"11",X"11",X"00",X"00",X"9F",X"99",X"00",X"00",X"99",X"F9",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"F0",X"90",X"00",X"00",X"9F",X"90",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"00",X"00",
		X"09",X"99",X"99",X"99",X"09",X"22",X"22",X"22",X"09",X"22",X"22",X"22",X"09",X"99",X"99",X"99",
		X"00",X"22",X"2C",X"99",X"00",X"22",X"22",X"22",X"00",X"9C",X"22",X"22",X"00",X"99",X"99",X"99",
		X"99",X"C9",X"22",X"22",X"22",X"9C",X"29",X"22",X"22",X"29",X"92",X"22",X"22",X"22",X"99",X"99",
		X"22",X"2C",X"99",X"99",X"22",X"2C",X"29",X"92",X"99",X"22",X"C2",X"22",X"09",X"99",X"99",X"29",
		X"09",X"29",X"99",X"99",X"09",X"C2",X"29",X"29",X"09",X"2C",X"22",X"22",X"09",X"2C",X"99",X"C2",
		X"09",X"99",X"99",X"C2",X"00",X"CC",X"29",X"99",X"00",X"CC",X"22",X"29",X"00",X"C2",X"2C",X"2C",
		X"00",X"C2",X"22",X"22",X"99",X"99",X"99",X"22",X"9C",X"99",X"92",X"C9",X"0C",X"22",X"2C",X"99",
		X"09",X"2C",X"22",X"33",X"09",X"2C",X"22",X"33",X"09",X"22",X"22",X"33",X"09",X"C2",X"22",X"33",
		X"99",X"99",X"99",X"FF",X"22",X"22",X"22",X"0F",X"22",X"22",X"22",X"00",X"99",X"99",X"99",X"00",
		X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"00",X"22",X"29",X"22",X"92",X"99",X"99",X"99",X"99",
		X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"29",X"22",X"32",X"22",X"2F",X"99",X"99",X"99",X"F0",
		X"00",X"00",X"FF",X"02",X"99",X"00",X"0F",X"0F",X"92",X"99",X"00",X"00",X"29",X"22",X"00",X"00",
		X"C2",X"22",X"20",X"FF",X"99",X"99",X"0F",X"00",X"22",X"92",X"2F",X"0F",X"29",X"29",X"00",X"0F",
		X"92",X"92",X"20",X"0F",X"99",X"92",X"00",X"00",X"CC",X"99",X"20",X"0F",X"22",X"22",X"0F",X"00",
		X"29",X"92",X"20",X"00",X"22",X"22",X"00",X"00",X"99",X"92",X"20",X"00",X"9C",X"99",X"00",X"00",
		X"CC",X"92",X"00",X"00",X"33",X"22",X"0F",X"0F",X"39",X"22",X"20",X"00",X"39",X"92",X"00",X"0F",
		X"00",X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"29",X"22",X"22",X"00",X"99",X"99",X"99",X"00",X"22",X"99",X"22",X"00",X"22",X"90",X"22",
		X"00",X"22",X"09",X"22",X"09",X"22",X"90",X"22",X"99",X"99",X"99",X"99",X"00",X"22",X"22",X"92",
		X"0C",X"22",X"92",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"29",X"29",X"00",X"99",X"29",X"33",
		X"09",X"99",X"92",X"22",X"09",X"92",X"29",X"29",X"09",X"C2",X"CC",X"22",X"00",X"C2",X"29",X"22",
		X"0F",X"C2",X"22",X"99",X"F9",X"C2",X"9F",X"00",X"09",X"99",X"FF",X"00",X"0F",X"29",X"0F",X"00",
		X"00",X"92",X"0F",X"00",X"0F",X"99",X"FF",X"00",X"F0",X"99",X"0F",X"00",X"0F",X"00",X"0F",X"00",
		X"F0",X"02",X"00",X"00",X"0F",X"F2",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"99",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"29",X"22",X"00",X"00",X"22",X"92",X"20",X"00",
		X"29",X"22",X"00",X"00",X"33",X"39",X"20",X"0F",X"22",X"22",X"00",X"00",X"29",X"92",X"20",X"00",
		X"22",X"22",X"00",X"00",X"99",X"22",X"20",X"0F",X"22",X"99",X"00",X"0F",X"29",X"22",X"20",X"00",
		X"29",X"22",X"00",X"0F",X"22",X"29",X"20",X"00",X"99",X"33",X"20",X"0F",X"39",X"29",X"20",X"00",
		X"93",X"22",X"00",X"F0",X"92",X"22",X"20",X"0F",X"29",X"99",X"0F",X"0F",X"99",X"F0",X"F2",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"0F",X"02",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"22",X"0F",
		X"00",X"00",X"20",X"0F",X"00",X"02",X"90",X"00",X"00",X"09",X"20",X"0F",X"00",X"99",X"0F",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"FF",X"00",
		X"09",X"99",X"99",X"99",X"09",X"22",X"22",X"22",X"09",X"22",X"22",X"22",X"09",X"99",X"99",X"99",
		X"00",X"22",X"2C",X"99",X"00",X"22",X"22",X"22",X"00",X"9C",X"22",X"22",X"00",X"99",X"99",X"99",
		X"99",X"C9",X"22",X"22",X"22",X"9C",X"29",X"22",X"22",X"29",X"92",X"22",X"22",X"22",X"99",X"99",
		X"22",X"2C",X"99",X"99",X"22",X"2C",X"29",X"92",X"99",X"22",X"C2",X"22",X"09",X"99",X"99",X"29",
		X"09",X"29",X"99",X"99",X"09",X"C2",X"29",X"29",X"09",X"2C",X"22",X"22",X"09",X"2C",X"99",X"C2",
		X"09",X"99",X"99",X"C2",X"00",X"CC",X"29",X"99",X"00",X"CC",X"22",X"29",X"00",X"C2",X"2C",X"2C",
		X"00",X"C2",X"22",X"22",X"99",X"99",X"99",X"22",X"9C",X"99",X"92",X"C9",X"0C",X"22",X"2C",X"99",
		X"09",X"2C",X"22",X"33",X"09",X"2C",X"22",X"33",X"09",X"22",X"22",X"33",X"09",X"C2",X"22",X"33",
		X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"FF",X"99",X"99",X"99",X"00",
		X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"00",X"22",X"29",X"22",X"92",X"99",X"99",X"99",X"99",
		X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"29",X"22",X"32",X"22",X"22",X"99",X"99",X"99",X"0F",
		X"00",X"00",X"00",X"F2",X"99",X"00",X"00",X"00",X"92",X"99",X"00",X"F0",X"29",X"22",X"00",X"00",
		X"C2",X"22",X"20",X"F0",X"99",X"99",X"00",X"00",X"22",X"92",X"20",X"00",X"29",X"29",X"20",X"F0",
		X"92",X"92",X"20",X"0F",X"99",X"92",X"92",X"FF",X"CC",X"99",X"22",X"00",X"22",X"22",X"29",X"00",
		X"29",X"92",X"29",X"0F",X"22",X"22",X"20",X"0F",X"99",X"92",X"20",X"0F",X"9C",X"99",X"29",X"00",
		X"CC",X"92",X"20",X"00",X"33",X"22",X"20",X"00",X"39",X"22",X"20",X"FF",X"39",X"92",X"99",X"FF",
		X"00",X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"29",X"22",X"22",X"00",X"99",X"99",X"99",X"00",X"22",X"99",X"22",X"00",X"22",X"90",X"22",
		X"00",X"22",X"09",X"22",X"09",X"22",X"90",X"22",X"99",X"99",X"99",X"99",X"00",X"22",X"22",X"92",
		X"0C",X"22",X"92",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"29",X"29",X"00",X"99",X"29",X"33",
		X"09",X"99",X"92",X"22",X"09",X"92",X"29",X"29",X"09",X"C2",X"CC",X"22",X"00",X"C2",X"29",X"22",
		X"00",X"C2",X"22",X"99",X"09",X"C2",X"92",X"00",X"09",X"99",X"02",X"00",X"00",X"29",X"02",X"00",
		X"00",X"92",X"FF",X"00",X"00",X"99",X"02",X"00",X"00",X"99",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"F2",X"00",X"00",X"00",X"F2",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"22",X"0F",X"22",X"22",X"20",X"F0",X"29",X"22",X"09",X"00",X"22",X"92",X"20",X"F0",
		X"29",X"22",X"F0",X"00",X"33",X"39",X"29",X"F0",X"22",X"22",X"20",X"0F",X"29",X"92",X"29",X"F0",
		X"22",X"22",X"90",X"00",X"99",X"22",X"2F",X"00",X"22",X"99",X"2F",X"00",X"29",X"22",X"20",X"00",
		X"29",X"22",X"F0",X"00",X"22",X"29",X"20",X"0F",X"99",X"33",X"20",X"00",X"39",X"29",X"20",X"0F",
		X"93",X"22",X"F0",X"00",X"92",X"22",X"2F",X"F0",X"29",X"99",X"00",X"00",X"99",X"00",X"F2",X"0F",
		X"00",X"00",X"0F",X"F0",X"00",X"00",X"02",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"22",X"0F",
		X"00",X"00",X"20",X"0F",X"00",X"02",X"90",X"0F",X"00",X"09",X"20",X"00",X"00",X"99",X"00",X"0F",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"3A",X"00",X"00",X"00",X"3E",X"AA",X"00",
		X"00",X"69",X"A9",X"AA",X"00",X"F9",X"9A",X"99",X"00",X"69",X"A9",X"99",X"00",X"99",X"99",X"99",
		X"0F",X"99",X"9A",X"A9",X"0F",X"F9",X"53",X"33",X"0F",X"F3",X"7A",X"F3",X"0F",X"FA",X"AA",X"FF",
		X"0F",X"F9",X"AA",X"55",X"0F",X"FF",X"AA",X"55",X"0F",X"FE",X"99",X"55",X"0F",X"FE",X"55",X"55",
		X"F5",X"EE",X"AA",X"55",X"F3",X"9E",X"AA",X"00",X"FF",X"9E",X"AA",X"FF",X"F0",X"A9",X"EA",X"55",
		X"F0",X"E9",X"AE",X"55",X"FF",X"5A",X"E5",X"55",X"FF",X"EE",X"EE",X"55",X"0F",X"E5",X"99",X"F5",
		X"F0",X"EE",X"99",X"FA",X"00",X"AA",X"99",X"AA",X"00",X"9F",X"99",X"EE",X"00",X"39",X"99",X"99",
		X"00",X"D0",X"D9",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"99",X"00",
		X"F9",X"9A",X"39",X"00",X"99",X"99",X"E3",X"00",X"0A",X"F9",X"99",X"0F",X"AA",X"99",X"99",X"0F",
		X"AA",X"77",X"99",X"90",X"AA",X"AA",X"59",X"90",X"AA",X"AA",X"75",X"40",X"AA",X"99",X"A7",X"90",
		X"AA",X"44",X"59",X"0F",X"AA",X"9A",X"79",X"0F",X"AA",X"A9",X"79",X"0F",X"AA",X"44",X"A9",X"0F",
		X"AA",X"9A",X"A9",X"0F",X"AA",X"44",X"A9",X"0F",X"AE",X"A9",X"A9",X"0F",X"EA",X"9A",X"E9",X"0F",
		X"EE",X"49",X"9F",X"F0",X"EE",X"A4",X"9F",X"F0",X"9E",X"EA",X"9F",X"F0",X"99",X"EE",X"99",X"F0",
		X"99",X"99",X"99",X"F0",X"D9",X"99",X"99",X"F0",X"09",X"99",X"9A",X"F0",X"00",X"3A",X"99",X"F0",
		X"00",X"93",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"05",X"55",X"99",X"00",
		X"05",X"AE",X"AE",X"0E",X"05",X"9A",X"9A",X"EE",X"59",X"99",X"A9",X"99",X"5F",X"A7",X"9A",X"9A",
		X"59",X"AA",X"99",X"AF",X"59",X"AA",X"A7",X"A9",X"5F",X"AA",X"EA",X"99",X"59",X"99",X"5E",X"A7",
		X"59",X"99",X"EE",X"EA",X"FF",X"39",X"5E",X"AE",X"99",X"99",X"EE",X"EA",X"99",X"9F",X"5E",X"AE",
		X"FF",X"EF",X"5E",X"EA",X"99",X"E9",X"E5",X"EE",X"99",X"E9",X"5E",X"AE",X"99",X"5E",X"E5",X"EE",
		X"33",X"9E",X"65",X"EE",X"06",X"A9",X"AA",X"E5",X"06",X"E9",X"DD",X"55",X"06",X"EA",X"FF",X"AA",
		X"00",X"EA",X"DD",X"DD",X"00",X"AE",X"AA",X"FF",X"00",X"0A",X"EE",X"DD",X"00",X"0E",X"00",X"AA",
		X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AE",X"00",X"00",X"00",
		X"EA",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"97",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"A9",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"EA",X"00",X"E5",
		X"96",X"AA",X"99",X"5E",X"96",X"EA",X"EA",X"99",X"96",X"A9",X"A9",X"A9",X"33",X"9A",X"FF",X"FF",
		X"99",X"99",X"A9",X"A9",X"99",X"79",X"99",X"99",X"9F",X"A9",X"A7",X"A7",X"FF",X"A9",X"EA",X"EA",
		X"99",X"9F",X"AE",X"AE",X"99",X"9F",X"EA",X"EA",X"FF",X"FF",X"AE",X"AE",X"99",X"F9",X"EE",X"EA",
		X"99",X"99",X"EE",X"AE",X"FF",X"F9",X"E5",X"EA",X"99",X"FF",X"5E",X"EE",X"99",X"9F",X"E5",X"EA",
		X"FF",X"9F",X"5E",X"5E",X"9F",X"E9",X"56",X"55",X"99",X"E9",X"AA",X"AA",X"99",X"99",X"DD",X"DD",
		X"33",X"AA",X"FF",X"FF",X"06",X"EA",X"DD",X"DD",X"06",X"EE",X"AA",X"AA",X"06",X"EA",X"EE",X"5E",
		X"00",X"AE",X"90",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"97",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"A9",X"00",X"00",X"00",X"DA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"99",X"00",
		X"09",X"5E",X"AA",X"9E",X"09",X"99",X"99",X"AA",X"99",X"99",X"33",X"EE",X"55",X"99",X"53",X"53",
		X"99",X"49",X"F0",X"33",X"55",X"44",X"5F",X"93",X"99",X"9A",X"55",X"39",X"55",X"91",X"FF",X"EB",
		X"99",X"44",X"FF",X"EE",X"55",X"99",X"FF",X"EA",X"99",X"94",X"FF",X"AE",X"59",X"1A",X"FF",X"EA",
		X"96",X"9A",X"55",X"EE",X"44",X"44",X"55",X"AE",X"9E",X"EE",X"55",X"EE",X"9F",X"99",X"F3",X"EE",
		X"9F",X"99",X"53",X"EE",X"99",X"99",X"39",X"B3",X"00",X"AA",X"95",X"99",X"00",X"AE",X"E5",X"99",
		X"00",X"99",X"AE",X"99",X"00",X"00",X"9A",X"99",X"00",X"00",X"09",X"3A",X"00",X"00",X"00",X"A9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"5A",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",
		X"5A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"A9",X"00",X"00",X"09",X"3A",X"00",X"00",X"9A",X"99",X"00",X"99",X"AE",X"99",
		X"00",X"EE",X"E5",X"99",X"00",X"EE",X"95",X"99",X"99",X"99",X"39",X"B3",X"9F",X"99",X"53",X"EE",
		X"9F",X"99",X"F3",X"EE",X"9E",X"EE",X"55",X"EE",X"44",X"44",X"55",X"AE",X"96",X"9A",X"55",X"EE",
		X"59",X"1A",X"FF",X"EA",X"99",X"94",X"FF",X"AE",X"55",X"99",X"FF",X"EA",X"99",X"44",X"FF",X"EE",
		X"55",X"91",X"FF",X"EB",X"99",X"9A",X"55",X"39",X"55",X"44",X"5F",X"93",X"99",X"49",X"F0",X"33",
		X"55",X"99",X"53",X"53",X"99",X"99",X"33",X"EE",X"09",X"99",X"99",X"AA",X"09",X"AE",X"AA",X"9E",
		X"00",X"AE",X"99",X"00",X"00",X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"33",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"90",X"90",X"99",X"00",X"09",X"02",X"92",X"09",X"99",X"99",X"22",
		X"99",X"99",X"99",X"22",X"21",X"A3",X"99",X"22",X"17",X"33",X"99",X"22",X"17",X"AA",X"29",X"22",
		X"31",X"3F",X"29",X"22",X"29",X"99",X"29",X"22",X"33",X"52",X"29",X"22",X"29",X"52",X"29",X"22",
		X"97",X"52",X"29",X"22",X"97",X"26",X"29",X"22",X"97",X"27",X"29",X"22",X"97",X"26",X"29",X"22",
		X"99",X"27",X"29",X"22",X"97",X"27",X"29",X"22",X"97",X"26",X"29",X"22",X"97",X"22",X"29",X"22",
		X"97",X"F2",X"29",X"22",X"29",X"F2",X"29",X"22",X"33",X"F9",X"29",X"22",X"39",X"92",X"29",X"22",
		X"21",X"3F",X"29",X"22",X"17",X"AA",X"29",X"22",X"17",X"33",X"09",X"22",X"21",X"A3",X"09",X"22",
		X"99",X"00",X"09",X"22",X"00",X"00",X"02",X"92",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"20",X"00",X"00",X"55",X"10",X"00",X"00",X"55",X"00",X"00",X"55",X"55",X"55",
		X"00",X"55",X"55",X"55",X"00",X"55",X"55",X"55",X"00",X"55",X"51",X"33",X"00",X"55",X"11",X"33",
		X"05",X"33",X"11",X"77",X"19",X"44",X"33",X"99",X"99",X"11",X"AB",X"33",X"55",X"13",X"BB",X"99",
		X"0F",X"55",X"BB",X"9D",X"00",X"53",X"9B",X"9D",X"00",X"33",X"B9",X"9D",X"01",X"33",X"B9",X"9D",
		X"01",X"53",X"B9",X"9D",X"00",X"53",X"B9",X"9D",X"00",X"F3",X"9B",X"9D",X"03",X"FF",X"BB",X"99",
		X"55",X"FF",X"BB",X"93",X"99",X"1F",X"AB",X"33",X"19",X"11",X"FF",X"FF",X"0F",X"55",X"11",X"11",
		X"00",X"55",X"11",X"55",X"00",X"55",X"51",X"55",X"00",X"55",X"55",X"FF",X"00",X"5F",X"55",X"FF",
		X"00",X"FF",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"10",X"00",X"00",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"09",X"99",X"00",X"00",
		X"99",X"9F",X"00",X"00",X"FF",X"F5",X"00",X"00",X"11",X"55",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"FF",X"00",X"00",X"99",X"9F",X"00",X"00",X"F9",X"99",X"00",X"00",
		X"0F",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"E9",X"99",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"E9",X"00",X"00",X"99",X"99",X"00",X"00",
		X"22",X"99",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"99",X"00",X"00",X"22",X"09",X"00",X"00",
		X"22",X"99",X"09",X"00",X"22",X"33",X"00",X"00",X"22",X"33",X"09",X"00",X"22",X"99",X"0F",X"00",
		X"22",X"99",X"9F",X"00",X"23",X"33",X"F9",X"00",X"22",X"33",X"F9",X"00",X"29",X"99",X"F9",X"00",
		X"22",X"99",X"99",X"00",X"22",X"99",X"9F",X"00",X"22",X"99",X"FF",X"00",X"22",X"29",X"99",X"00",
		X"99",X"92",X"99",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"9F",X"00",
		X"22",X"22",X"9F",X"00",X"22",X"22",X"9F",X"00",X"99",X"99",X"9F",X"00",X"22",X"22",X"FF",X"00",
		X"22",X"22",X"F9",X"00",X"22",X"22",X"F0",X"00",X"22",X"22",X"99",X"00",X"22",X"22",X"90",X"00",
		X"11",X"11",X"90",X"00",X"11",X"11",X"99",X"00",X"11",X"11",X"F0",X"00",X"11",X"11",X"F9",X"00",
		X"11",X"11",X"FF",X"00",X"11",X"11",X"9F",X"00",X"11",X"21",X"9F",X"00",X"12",X"22",X"9F",X"00",
		X"11",X"11",X"9F",X"00",X"11",X"91",X"99",X"00",X"11",X"11",X"99",X"00",X"11",X"11",X"99",X"00",
		X"11",X"19",X"99",X"00",X"11",X"99",X"FF",X"00",X"11",X"99",X"9F",X"00",X"22",X"99",X"99",X"00",
		X"19",X"99",X"F9",X"00",X"11",X"33",X"F9",X"00",X"13",X"33",X"F9",X"00",X"11",X"99",X"9F",X"00",
		X"11",X"99",X"0F",X"00",X"11",X"33",X"09",X"00",X"22",X"33",X"00",X"00",X"11",X"99",X"09",X"00",
		X"11",X"09",X"00",X"00",X"11",X"99",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"99",X"00",X"00",
		X"99",X"99",X"00",X"00",X"EE",X"E9",X"00",X"00",X"EE",X"90",X"00",X"00",X"E9",X"99",X"00",X"00",
		X"09",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"15",X"00",X"00",X"55",X"11",X"50",X"00",X"95",X"11",X"55",X"00",
		X"91",X"11",X"55",X"00",X"99",X"51",X"55",X"00",X"19",X"55",X"55",X"00",X"11",X"55",X"55",X"00",
		X"11",X"53",X"55",X"00",X"51",X"33",X"55",X"00",X"51",X"55",X"11",X"00",X"55",X"F5",X"11",X"50",
		X"55",X"F5",X"11",X"11",X"F5",X"5F",X"11",X"99",X"F5",X"F5",X"11",X"99",X"F5",X"F9",X"F1",X"99",
		X"F5",X"F9",X"BF",X"99",X"FF",X"F9",X"BB",X"09",X"0F",X"F9",X"9B",X"09",X"0F",X"F9",X"99",X"00",
		X"0F",X"FF",X"19",X"F0",X"00",X"1F",X"11",X"50",X"00",X"11",X"59",X"5F",X"00",X"11",X"99",X"5F",
		X"00",X"11",X"99",X"55",X"00",X"11",X"9D",X"25",X"00",X"11",X"9D",X"15",X"00",X"19",X"09",X"12",
		X"11",X"20",X"F9",X"99",X"11",X"11",X"FF",X"99",X"19",X"11",X"FF",X"FF",X"19",X"55",X"F9",X"0F",
		X"19",X"55",X"99",X"00",X"09",X"FF",X"9F",X"99",X"09",X"00",X"F9",X"99",X"00",X"90",X"39",X"FF",
		X"00",X"09",X"3F",X"1F",X"00",X"90",X"13",X"11",X"00",X"00",X"11",X"31",X"00",X"00",X"F1",X"31",
		X"00",X"00",X"F1",X"F3",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"F9",X"F9",
		X"00",X"00",X"F9",X"99",X"00",X"00",X"F9",X"09",X"00",X"00",X"F9",X"90",X"00",X"00",X"F9",X"09",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"6F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"09",X"00",X"09",X"33",X"00",X"00",X"09",X"53",X"99",X"00",X"0F",X"55",X"33",X"90",
		X"01",X"55",X"F3",X"09",X"11",X"11",X"5F",X"90",X"1F",X"11",X"5F",X"99",X"1F",X"11",X"55",X"33",
		X"01",X"55",X"55",X"FF",X"91",X"55",X"15",X"11",X"99",X"55",X"11",X"11",X"19",X"55",X"11",X"11",
		X"51",X"55",X"F1",X"11",X"55",X"F5",X"5F",X"19",X"55",X"FF",X"9B",X"99",X"F5",X"FF",X"BB",X"99",
		X"0F",X"FF",X"BB",X"95",X"0F",X"1F",X"B9",X"11",X"00",X"11",X"B9",X"B1",X"00",X"11",X"99",X"99",
		X"00",X"51",X"B9",X"99",X"00",X"55",X"BB",X"9D",X"00",X"5F",X"FB",X"DD",X"00",X"55",X"11",X"DF",
		X"00",X"55",X"11",X"DF",X"00",X"55",X"11",X"FF",X"00",X"F5",X"11",X"99",X"00",X"FF",X"11",X"11",
		X"00",X"FF",X"11",X"51",X"00",X"0F",X"11",X"5F",X"00",X"00",X"11",X"FF",X"00",X"00",X"11",X"FF",
		X"55",X"F5",X"90",X"00",X"11",X"5F",X"90",X"00",X"11",X"55",X"90",X"00",X"11",X"51",X"99",X"00",
		X"95",X"11",X"90",X"00",X"5F",X"11",X"90",X"00",X"55",X"11",X"09",X"00",X"FF",X"11",X"90",X"00",
		X"F9",X"11",X"39",X"00",X"F9",X"BF",X"33",X"00",X"F9",X"9B",X"F3",X"00",X"F9",X"29",X"F3",X"00",
		X"F9",X"22",X"59",X"00",X"FB",X"22",X"5F",X"90",X"1F",X"51",X"5F",X"F9",X"11",X"51",X"9F",X"FF",
		X"11",X"99",X"19",X"00",X"11",X"99",X"F1",X"99",X"51",X"1F",X"F8",X"FF",X"52",X"11",X"F8",X"99",
		X"55",X"51",X"88",X"FF",X"55",X"55",X"8F",X"FF",X"F5",X"5F",X"19",X"11",X"F5",X"FF",X"11",X"55",
		X"FF",X"0F",X"F1",X"55",X"FF",X"00",X"FF",X"55",X"0F",X"00",X"F9",X"5F",X"00",X"00",X"F9",X"9F",
		X"00",X"00",X"F9",X"F3",X"00",X"00",X"FF",X"F3",X"00",X"00",X"9F",X"0F",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",
		X"99",X"CC",X"99",X"99",X"99",X"EB",X"99",X"99",X"59",X"AA",X"CC",X"99",X"59",X"AC",X"00",X"99",
		X"C5",X"AB",X"EB",X"CC",X"C5",X"EE",X"AA",X"9B",X"C5",X"BE",X"BE",X"C9",X"CF",X"BB",X"EB",X"BC",
		X"CF",X"BB",X"BB",X"BB",X"CF",X"EE",X"5B",X"9B",X"C5",X"F5",X"BB",X"CB",X"CF",X"BB",X"BB",X"B9",
		X"5E",X"BB",X"BB",X"9A",X"99",X"BB",X"5B",X"9A",X"65",X"BB",X"B5",X"9A",X"65",X"BB",X"5B",X"9A",
		X"65",X"96",X"BF",X"99",X"CB",X"BB",X"FB",X"9B",X"0C",X"CC",X"BB",X"BB",X"00",X"BB",X"6F",X"B9",
		X"0C",X"9B",X"BF",X"CC",X"00",X"09",X"CB",X"BC",X"00",X"00",X"9C",X"BB",X"00",X"00",X"09",X"BB",
		X"00",X"00",X"00",X"CC",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",
		X"00",X"00",X"99",X"9C",X"00",X"90",X"99",X"BB",X"00",X"99",X"9C",X"99",X"00",X"99",X"CB",X"BC",
		X"00",X"9B",X"AA",X"CC",X"09",X"BB",X"BA",X"B9",X"0C",X"CC",X"AB",X"BB",X"CB",X"AA",X"BB",X"9B",
		X"65",X"9A",X"BB",X"99",X"65",X"BB",X"BB",X"9A",X"65",X"AB",X"BB",X"9A",X"99",X"BB",X"BB",X"9A",
		X"5E",X"BB",X"BB",X"9A",X"CF",X"BB",X"BB",X"B9",X"C5",X"EE",X"B5",X"CB",X"CF",X"F5",X"5B",X"9B",
		X"CF",X"BB",X"BF",X"5B",X"CF",X"BB",X"5B",X"BC",X"C5",X"BE",X"B5",X"C9",X"C5",X"EE",X"FA",X"9B",
		X"C5",X"AB",X"EB",X"CC",X"59",X"BB",X"00",X"AA",X"00",X"6B",X"CC",X"00",X"00",X"EB",X"AA",X"00",
		X"00",X"CC",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"99",X"00",X"D0",X"D9",X"99",
		X"00",X"39",X"99",X"99",X"00",X"9F",X"99",X"EE",X"00",X"AA",X"99",X"AA",X"F0",X"EE",X"99",X"FA",
		X"0F",X"E5",X"99",X"F5",X"FF",X"EE",X"EE",X"55",X"FF",X"5A",X"E5",X"55",X"F0",X"E9",X"AE",X"55",
		X"F0",X"A9",X"EA",X"55",X"FF",X"9E",X"AA",X"FF",X"F3",X"9E",X"AA",X"00",X"F5",X"EE",X"AA",X"55",
		X"0F",X"FE",X"55",X"55",X"0F",X"FE",X"99",X"55",X"0F",X"FF",X"AA",X"55",X"0F",X"F9",X"AA",X"55",
		X"0F",X"FA",X"AA",X"FF",X"0F",X"F3",X"7A",X"F3",X"0F",X"F9",X"53",X"33",X"0F",X"99",X"9A",X"A9",
		X"00",X"99",X"99",X"99",X"00",X"69",X"A9",X"99",X"00",X"F9",X"9A",X"99",X"00",X"69",X"A9",X"AA",
		X"00",X"3E",X"AA",X"00",X"00",X"3A",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"93",X"99",X"00",
		X"00",X"3A",X"99",X"F0",X"09",X"99",X"9A",X"F0",X"D9",X"99",X"99",X"F0",X"99",X"99",X"99",X"F0",
		X"99",X"EE",X"99",X"F0",X"9E",X"EA",X"9F",X"F0",X"EE",X"A4",X"9F",X"F0",X"EE",X"49",X"9F",X"F0",
		X"EA",X"9A",X"E9",X"0F",X"AE",X"A9",X"A9",X"0F",X"AA",X"44",X"A9",X"0F",X"AA",X"9A",X"A9",X"0F",
		X"AA",X"44",X"A9",X"0F",X"AA",X"A9",X"79",X"0F",X"AA",X"9A",X"79",X"0F",X"AA",X"44",X"59",X"0F",
		X"AA",X"99",X"A7",X"90",X"AA",X"AA",X"75",X"40",X"AA",X"AA",X"59",X"90",X"AA",X"77",X"99",X"90",
		X"AA",X"99",X"99",X"0F",X"0A",X"F9",X"99",X"0F",X"99",X"99",X"E3",X"00",X"F9",X"9A",X"39",X"00",
		X"99",X"99",X"99",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"22",X"09",X"90",
		X"9F",X"2D",X"99",X"90",X"96",X"11",X"22",X"29",X"92",X"11",X"22",X"22",X"92",X"71",X"99",X"22",
		X"F2",X"11",X"33",X"22",X"52",X"11",X"11",X"99",X"52",X"11",X"DD",X"33",X"52",X"D1",X"77",X"11",
		X"52",X"41",X"77",X"DA",X"52",X"41",X"77",X"7D",X"52",X"41",X"57",X"7D",X"52",X"71",X"77",X"77",
		X"2D",X"59",X"77",X"51",X"2E",X"19",X"57",X"71",X"27",X"1F",X"77",X"71",X"67",X"19",X"57",X"51",
		X"F2",X"19",X"F7",X"71",X"22",X"11",X"11",X"51",X"90",X"77",X"33",X"71",X"00",X"22",X"99",X"11",
		X"00",X"22",X"29",X"91",X"00",X"90",X"52",X"99",X"00",X"00",X"22",X"22",X"00",X"00",X"02",X"52",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",X"1F",X"00",X"00",X"00",
		X"1F",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"22",
		X"00",X"00",X"99",X"22",X"00",X"99",X"22",X"22",X"00",X"99",X"22",X"99",X"00",X"22",X"29",X"91",
		X"90",X"22",X"99",X"11",X"99",X"77",X"33",X"77",X"22",X"11",X"11",X"57",X"F2",X"19",X"D7",X"77",
		X"67",X"19",X"77",X"71",X"27",X"19",X"77",X"71",X"2E",X"19",X"77",X"71",X"2D",X"59",X"77",X"51",
		X"52",X"71",X"77",X"77",X"52",X"41",X"57",X"7D",X"52",X"41",X"77",X"5D",X"52",X"41",X"77",X"DA",
		X"52",X"D1",X"55",X"11",X"52",X"11",X"55",X"33",X"52",X"11",X"11",X"99",X"F2",X"11",X"33",X"22",
		X"92",X"71",X"99",X"22",X"92",X"11",X"22",X"55",X"96",X"11",X"52",X"20",X"9F",X"2D",X"00",X"00",
		X"99",X"22",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"77",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"15",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"95",X"00",X"00",X"93",X"55",X"00",X"00",X"55",X"50",X"00",X"00",X"55",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"5F",X"90",X"00",
		X"00",X"5F",X"59",X"00",X"00",X"0F",X"55",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"9A",X"9A",X"00",X"AB",X"AB",X"AB",X"00",X"BD",X"BD",X"BD",X"00",X"BB",X"BB",X"BB",
		X"00",X"5B",X"5B",X"5B",X"00",X"BA",X"BA",X"BA",X"00",X"DD",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"DD",X"EE",X"55",X"00",X"99",X"B5",X"99",X"00",X"DD",X"5B",X"EE",X"09",X"99",X"B5",X"99",
		X"9D",X"DD",X"99",X"99",X"99",X"99",X"F5",X"9A",X"DD",X"D9",X"5F",X"99",X"99",X"9E",X"FF",X"9A",
		X"AA",X"9A",X"5F",X"99",X"AB",X"A5",X"FF",X"9A",X"BA",X"BA",X"5F",X"99",X"0B",X"AB",X"55",X"9A",
		X"0A",X"BA",X"5B",X"99",X"00",X"AB",X"B5",X"FF",X"00",X"BA",X"5B",X"99",X"00",X"AB",X"F5",X"F5",
		X"00",X"BA",X"99",X"99",X"00",X"AB",X"55",X"99",X"00",X"99",X"99",X"99",X"00",X"BA",X"BA",X"BA",
		X"00",X"AB",X"AB",X"AB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"AB",X"AB",X"AB",
		X"99",X"99",X"99",X"00",X"AB",X"AB",X"AB",X"00",X"BD",X"BD",X"BD",X"00",X"BB",X"BB",X"BB",X"00",
		X"5B",X"5B",X"5B",X"00",X"BA",X"BA",X"BA",X"00",X"99",X"DD",X"DD",X"00",X"99",X"DD",X"DD",X"00",
		X"99",X"BB",X"BB",X"00",X"9E",X"DD",X"DD",X"00",X"EA",X"BB",X"BB",X"00",X"AE",X"DD",X"DD",X"00",
		X"EA",X"BB",X"BB",X"00",X"AE",X"BD",X"DB",X"00",X"AA",X"BB",X"BB",X"00",X"A9",X"BB",X"BB",X"00",
		X"9A",X"BB",X"AB",X"00",X"AA",X"BB",X"BB",X"00",X"9A",X"AB",X"AB",X"00",X"A9",X"BB",X"BB",X"00",
		X"99",X"AA",X"AA",X"00",X"99",X"BB",X"BB",X"00",X"99",X"AA",X"AA",X"00",X"59",X"B9",X"B9",X"00",
		X"55",X"AA",X"AA",X"00",X"55",X"B9",X"99",X"00",X"99",X"99",X"99",X"00",X"AB",X"AB",X"AB",X"00",
		X"BA",X"BA",X"BA",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"AB",X"AB",X"AB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"B0",
		X"0B",X"FB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"0B",X"00",X"BB",X"BB",
		X"0B",X"00",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"BB",X"0B",X"0B",X"BB",X"BB",X"00",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",
		X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"FB",X"00",X"BB",X"00",X"BB",X"00",X"BB",
		X"00",X"BB",X"00",X"FB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",
		X"0B",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"BB",X"0B",X"BF",X"FF",X"BB",X"0B",X"FB",X"BB",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"FB",X"00",X"0B",X"BB",X"BF",X"B0",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"FF",X"00",X"BB",X"BB",X"BB",X"0B",X"00",X"BB",X"BB",
		X"0B",X"00",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"BB",X"0B",X"0B",X"BB",X"BB",X"00",
		X"0B",X"FB",X"BB",X"BB",X"0B",X"FB",X"BB",X"FB",X"0B",X"FB",X"BB",X"FF",X"0B",X"FB",X"BB",X"FF",
		X"0B",X"FB",X"00",X"BF",X"0B",X"FB",X"00",X"BF",X"0B",X"FB",X"00",X"BF",X"0B",X"FB",X"00",X"BF",
		X"0B",X"FB",X"00",X"BF",X"0B",X"FB",X"00",X"BF",X"0B",X"FB",X"00",X"BF",X"0B",X"FB",X"00",X"BF",
		X"0B",X"FF",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",
		X"00",X"BB",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",
		X"0B",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"FF",X"FF",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"BB",X"FF",X"0B",X"BB",X"BB",X"BF",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"FB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"FF",X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"FF",X"B0",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"0B",X"00",X"BB",X"BB",
		X"0B",X"00",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"BB",X"0B",X"0B",X"BB",X"FF",X"00",
		X"0B",X"BB",X"FB",X"BB",X"0B",X"BB",X"FF",X"BB",X"0B",X"BB",X"FF",X"BB",X"0B",X"BB",X"BB",X"BB",
		X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"FB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"FB",X"00",X"FB",X"00",X"BB",X"00",X"FB",X"00",X"BB",X"00",X"FF",X"00",X"BB",X"00",X"BF",
		X"00",X"BB",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",
		X"0B",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BF",X"FF",X"BB",
		X"00",X"FF",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"FB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"B0",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"FB",X"BB",X"BB",
		X"0B",X"FF",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"00",X"BB",X"FF",X"BB",X"0B",X"00",X"BB",X"BB",
		X"0B",X"00",X"00",X"FB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"BB",X"0B",X"0B",X"BB",X"BB",X"00",
		X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"BB",X"BB",
		X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",X"00",X"BB",
		X"0B",X"BB",X"00",X"BB",X"00",X"FB",X"00",X"BB",X"00",X"FF",X"00",X"FB",X"00",X"FB",X"00",X"FB",
		X"00",X"BB",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"0B",
		X"0B",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BB",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"BB",
		X"00",X"BB",X"FB",X"BB",X"0B",X"BF",X"FF",X"BB",X"0B",X"FF",X"BB",X"BB",X"0B",X"FB",X"00",X"BB",
		X"0B",X"B0",X"00",X"FB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",
		X"0B",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"00",X"01",X"11",X"11",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"11",X"01",X"11",X"01",X"11",X"01",X"11",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"01",X"11",X"01",X"11",X"01",X"11",X"01",X"11",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"01",X"01",X"11",X"11",X"11",X"00",X"00",X"01",X"11",
		X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"01",X"11",X"00",
		X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"00",X"01",X"11",X"11",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"11",X"01",X"00",X"01",X"11",X"01",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"11",X"01",X"01",X"01",X"11",X"01",X"11",
		X"01",X"00",X"01",X"11",X"01",X"00",X"01",X"10",X"01",X"00",X"01",X"00",X"01",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"01",X"11",X"01",X"11",X"01",X"11",
		X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"11",X"11",X"11",X"01",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",
		X"01",X"00",X"11",X"00",X"01",X"00",X"11",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"E6",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E6",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"E6",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"E0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",X"09",X"09",X"00",X"99",X"99",X"99",
		X"09",X"55",X"99",X"5F",X"EE",X"EE",X"EE",X"EE",X"EB",X"BB",X"BB",X"BB",X"E4",X"42",X"99",X"11",
		X"F7",X"77",X"99",X"99",X"F3",X"55",X"55",X"99",X"F5",X"55",X"FF",X"55",X"55",X"55",X"FF",X"F5",
		X"F5",X"55",X"FF",X"59",X"F5",X"B5",X"FF",X"59",X"F5",X"55",X"FF",X"59",X"F5",X"55",X"FF",X"59",
		X"F5",X"55",X"FF",X"59",X"F5",X"55",X"FF",X"59",X"F5",X"FF",X"FF",X"59",X"F5",X"55",X"FF",X"59",
		X"55",X"55",X"FF",X"F5",X"F5",X"55",X"FF",X"55",X"F3",X"55",X"55",X"99",X"FF",X"77",X"99",X"99",
		X"FF",X"42",X"99",X"11",X"EF",X"BB",X"BB",X"BB",X"EE",X"FF",X"FF",X"FF",X"00",X"55",X"00",X"5F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9B",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"09",X"00",X"00",
		X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"9B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
