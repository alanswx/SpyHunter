library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity spy_hunter_sp_bits_3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(14 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of spy_hunter_sp_bits_3 is
	type rom is array(0 to  32767) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"17",X"00",
		X"00",X"00",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"49",
		X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"00",X"00",X"00",X"23",X"00",X"00",X"00",X"17",X"00",
		X"00",X"00",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"99",X"00",X"00",X"BA",X"AA",X"AA",X"00",X"EB",X"AA",X"EE",X"0B",X"BB",X"AA",X"EB",
		X"EB",X"99",X"AA",X"BE",X"BB",X"99",X"99",X"EB",X"BB",X"99",X"BB",X"BE",X"BB",X"9B",X"BB",X"BB",
		X"BB",X"BB",X"55",X"5B",X"BA",X"B5",X"55",X"55",X"BA",X"B5",X"FF",X"55",X"55",X"55",X"AF",X"F5",
		X"BA",X"B5",X"FF",X"55",X"BA",X"B5",X"55",X"55",X"BB",X"BB",X"65",X"5B",X"BB",X"9B",X"BB",X"BB",
		X"BB",X"99",X"BB",X"BE",X"BB",X"99",X"99",X"EB",X"EB",X"99",X"AA",X"BE",X"0B",X"BB",X"AA",X"EB",
		X"00",X"EB",X"AA",X"EE",X"00",X"BA",X"AA",X"AA",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"EE",X"AA",X"00",X"00",
		X"AB",X"EE",X"E0",X"00",X"55",X"B5",X"EA",X"00",X"55",X"55",X"B5",X"AA",X"FF",X"FF",X"FF",X"5B",
		X"55",X"55",X"B5",X"AA",X"55",X"B5",X"EA",X"00",X"AB",X"EE",X"E0",X"00",X"EE",X"AA",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"99",X"00",X"99",X"BA",X"09",X"00",X"09",X"BB",X"09",X"00",X"00",X"AB",X"99",X"00",
		X"0B",X"99",X"90",X"00",X"BB",X"AA",X"99",X"99",X"BB",X"AA",X"A9",X"99",X"BB",X"99",X"AA",X"09",
		X"BB",X"9B",X"AA",X"09",X"BB",X"BB",X"AA",X"99",X"BB",X"B5",X"EA",X"99",X"BB",X"55",X"BE",X"AA",
		X"BB",X"5F",X"BB",X"AA",X"BB",X"55",X"5B",X"EB",X"BB",X"55",X"55",X"BE",X"AB",X"B5",X"55",X"EB",
		X"0A",X"BB",X"F5",X"BE",X"0A",X"BB",X"FF",X"BB",X"00",X"BB",X"55",X"BB",X"00",X"BB",X"55",X"BB",
		X"00",X"BA",X"B5",X"55",X"00",X"AA",X"BB",X"55",X"00",X"9A",X"9B",X"FF",X"00",X"99",X"9B",X"5F",
		X"00",X"90",X"9B",X"55",X"00",X"00",X"EB",X"B5",X"00",X"90",X"EB",X"BB",X"00",X"99",X"99",X"BB",
		X"00",X"09",X"A9",X"EB",X"00",X"00",X"09",X"AA",X"00",X"00",X"99",X"AA",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"BA",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"5B",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"BB",X"AE",X"00",X"00",
		X"AB",X"BB",X"00",X"00",X"AA",X"5B",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"FA",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"90",X"00",X"BA",X"9B",X"99",X"00",X"AA",X"A9",X"99",X"00",
		X"AA",X"A9",X"09",X"00",X"AA",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",X"AA",X"99",X"00",X"00",
		X"AA",X"BB",X"00",X"00",X"AA",X"BB",X"00",X"00",X"FA",X"BB",X"90",X"00",X"99",X"5B",X"90",X"00",
		X"99",X"55",X"99",X"00",X"99",X"55",X"99",X"00",X"9B",X"A5",X"99",X"00",X"BB",X"A5",X"99",X"00",
		X"BB",X"FF",X"99",X"90",X"BB",X"FF",X"9B",X"90",X"BA",X"5F",X"BE",X"00",X"AA",X"5F",X"EB",X"00",
		X"9A",X"55",X"BE",X"00",X"0A",X"B5",X"EB",X"00",X"09",X"B5",X"BE",X"00",X"00",X"BB",X"EB",X"00",
		X"00",X"BB",X"BE",X"00",X"00",X"EB",X"EB",X"00",X"00",X"BE",X"BE",X"00",X"90",X"EB",X"BB",X"00",
		X"90",X"BE",X"BC",X"00",X"99",X"AB",X"BB",X"00",X"09",X"AA",X"5B",X"00",X"09",X"00",X"5B",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"B5",X"00",
		X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AB",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"A0",
		X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"BA",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",
		X"00",X"90",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"9B",X"90",X"00",X"00",X"9B",X"9E",X"00",
		X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"AA",X"AB",X"00",X"00",X"FA",X"AA",X"00",
		X"00",X"AA",X"AA",X"00",X"00",X"FA",X"AA",X"00",X"00",X"FA",X"AA",X"00",X"00",X"9F",X"9A",X"00",
		X"00",X"9B",X"99",X"00",X"00",X"BB",X"B9",X"00",X"90",X"BB",X"BB",X"90",X"90",X"B5",X"BB",X"90",
		X"99",X"BB",X"BB",X"90",X"90",X"B5",X"B9",X"90",X"90",X"B5",X"B9",X"90",X"90",X"BB",X"BB",X"90",
		X"90",X"B5",X"B9",X"90",X"90",X"BB",X"B9",X"90",X"90",X"B5",X"B9",X"90",X"90",X"B5",X"B9",X"90",
		X"90",X"BB",X"B9",X"90",X"90",X"B5",X"B9",X"90",X"99",X"B5",X"B9",X"90",X"99",X"BB",X"BB",X"90",
		X"99",X"B5",X"BB",X"90",X"90",X"BB",X"BE",X"90",X"90",X"BB",X"BB",X"90",X"90",X"BB",X"BE",X"90",
		X"00",X"EB",X"EB",X"00",X"00",X"BB",X"BE",X"00",X"00",X"EB",X"EB",X"00",X"00",X"BE",X"BE",X"00",
		X"00",X"EB",X"EA",X"00",X"00",X"EB",X"EA",X"00",X"00",X"AB",X"A0",X"00",X"00",X"AE",X"A0",X"00",
		X"00",X"AB",X"A0",X"00",X"00",X"AB",X"A0",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"0F",X"53",X"00",X"00",X"F0",X"03",
		X"00",X"00",X"50",X"FF",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"03",X"00",X"05",X"00",X"0F",
		X"00",X"50",X"00",X"F0",X"00",X"55",X"00",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"50",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"50",X"00",X"0F",X"0F",X"00",X"00",X"F0",
		X"0F",X"05",X"00",X"00",X"0F",X"5F",X"00",X"05",X"0F",X"5F",X"00",X"F0",X"FF",X"5F",X"50",X"00",
		X"FF",X"53",X"00",X"00",X"FF",X"F0",X"33",X"00",X"FF",X"F0",X"00",X"35",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F5",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"F5",X"00",
		X"00",X"50",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"0F",X"05",X"00",X"00",X"3F",X"00",X"00",
		X"00",X"0F",X"3F",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F0",X"F0",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"50",X"05",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"05",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"05",X"00",X"00",X"03",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"39",
		X"FF",X"00",X"00",X"30",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"90",X"90",X"00",X"00",X"59",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"44",X"00",X"00",X"44",X"66",X"00",X"00",X"61",X"1F",X"00",X"0F",X"66",X"FF",
		X"00",X"00",X"44",X"66",X"00",X"00",X"06",X"44",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"19",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"06",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"FA",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"A0",X"05",X"00",X"00",X"A0",X"05",X"00",X"00",X"A0",X"50",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"A0",X"E0",X"55",X"00",X"5A",X"E0",X"55",X"00",
		X"5A",X"EF",X"5A",X"00",X"5A",X"EF",X"AE",X"00",X"5A",X"EF",X"AE",X"00",X"F0",X"A5",X"AE",X"00",
		X"00",X"AF",X"AE",X"00",X"00",X"A5",X"AE",X"00",X"0F",X"A5",X"AE",X"00",X"0F",X"5E",X"AE",X"00",
		X"0F",X"55",X"AE",X"00",X"00",X"55",X"AE",X"00",X"00",X"55",X"AE",X"00",X"00",X"5E",X"AA",X"00",
		X"00",X"5E",X"5A",X"00",X"00",X"55",X"5A",X"00",X"00",X"F5",X"55",X"00",X"00",X"55",X"55",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"00",
		X"99",X"09",X"99",X"00",X"90",X"09",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"90",X"00",
		X"99",X"99",X"00",X"00",X"90",X"99",X"00",X"00",X"00",X"D9",X"90",X"00",X"99",X"DD",X"90",X"00",
		X"90",X"99",X"99",X"00",X"99",X"09",X"99",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"09",X"99",X"00",X"00",X"09",X"99",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"99",X"99",X"09",X"00",X"09",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"90",X"00",X"99",X"99",X"00",X"99",X"99",X"99",X"00",
		X"9D",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"53",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"55",X"00",X"00",X"05",X"55",X"00",X"00",X"55",X"55",X"00",X"00",X"F5",X"55",X"00",
		X"00",X"0F",X"55",X"00",X"00",X"0F",X"55",X"00",X"00",X"3F",X"30",X"00",X"33",X"55",X"53",X"00",
		X"EE",X"35",X"55",X"00",X"5E",X"53",X"55",X"00",X"55",X"55",X"33",X"00",X"00",X"F5",X"E3",X"00",
		X"00",X"FF",X"55",X"00",X"35",X"00",X"5E",X"00",X"EE",X"05",X"E5",X"00",X"5E",X"55",X"55",X"00",
		X"F5",X"50",X"F5",X"00",X"F5",X"5F",X"55",X"00",X"05",X"FF",X"0F",X"00",X"00",X"5F",X"F5",X"00",
		X"00",X"55",X"F5",X"00",X"00",X"55",X"05",X"00",X"00",X"F5",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"55",X"05",X"00",X"00",X"50",X"F5",X"00",X"00",X"55",X"F5",X"00",
		X"00",X"E5",X"FF",X"30",X"00",X"5E",X"5F",X"30",X"00",X"55",X"55",X"E3",X"00",X"55",X"55",X"50",
		X"00",X"55",X"F5",X"00",X"00",X"5E",X"55",X"00",X"00",X"55",X"F5",X"00",X"00",X"55",X"55",X"00",
		X"00",X"5F",X"F5",X"30",X"00",X"F5",X"E5",X"E3",X"00",X"F5",X"5E",X"5E",X"00",X"5F",X"55",X"5E",
		X"00",X"F5",X"F5",X"5E",X"00",X"5F",X"55",X"30",X"00",X"5F",X"55",X"30",X"00",X"55",X"55",X"00",
		X"00",X"55",X"55",X"00",X"0F",X"55",X"5F",X"00",X"00",X"55",X"F5",X"00",X"00",X"55",X"F5",X"00",
		X"00",X"5F",X"FF",X"00",X"00",X"F5",X"F5",X"00",X"00",X"5F",X"0F",X"00",X"00",X"EF",X"00",X"00",
		X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F9",X"00",X"00",X"0E",X"EF",X"00",X"00",X"0F",X"BE",X"09",X"00",X"5F",X"4B",X"99",X"00",
		X"9F",X"4B",X"99",X"00",X"55",X"74",X"EE",X"00",X"F5",X"57",X"BB",X"90",X"F5",X"55",X"99",X"99",
		X"F5",X"55",X"99",X"55",X"F5",X"55",X"55",X"EE",X"F5",X"55",X"FF",X"BB",X"55",X"59",X"F5",X"15",
		X"99",X"59",X"FF",X"99",X"F9",X"59",X"FF",X"99",X"5F",X"93",X"FF",X"5B",X"55",X"93",X"FF",X"59",
		X"35",X"93",X"FF",X"99",X"73",X"93",X"FF",X"99",X"75",X"33",X"FF",X"99",X"47",X"93",X"FF",X"99",
		X"B4",X"99",X"FF",X"99",X"FF",X"93",X"FF",X"99",X"5F",X"55",X"FF",X"99",X"05",X"BF",X"FF",X"99",
		X"00",X"FB",X"FF",X"99",X"00",X"FF",X"FF",X"E3",X"00",X"00",X"9F",X"55",X"00",X"00",X"BB",X"55",
		X"00",X"00",X"FE",X"5F",X"00",X"00",X"00",X"54",X"00",X"00",X"05",X"BB",X"00",X"00",X"00",X"FB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",
		X"EA",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"43",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",X"A5",X"00",X"00",X"00",
		X"A9",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"54",X"00",X"00",X"02",X"55",X"00",X"00",X"92",X"55",X"90",X"00",X"99",X"F5",X"00",X"00",
		X"F3",X"FF",X"90",X"00",X"53",X"5F",X"99",X"00",X"75",X"5F",X"90",X"00",X"55",X"55",X"99",X"00",
		X"55",X"55",X"99",X"00",X"75",X"B5",X"A9",X"00",X"75",X"B5",X"A9",X"00",X"75",X"B5",X"A9",X"00",
		X"77",X"B5",X"EA",X"00",X"47",X"55",X"EA",X"00",X"47",X"55",X"EA",X"00",X"E7",X"99",X"EA",X"00",
		X"E4",X"99",X"EE",X"00",X"E4",X"99",X"9E",X"00",X"AE",X"99",X"9E",X"00",X"AE",X"99",X"9E",X"00",
		X"AE",X"99",X"9E",X"00",X"0A",X"9F",X"99",X"00",X"0A",X"FF",X"99",X"00",X"0A",X"FF",X"99",X"00",
		X"0A",X"FF",X"99",X"00",X"00",X"FF",X"59",X"90",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"F5",X"90",
		X"00",X"FF",X"95",X"00",X"00",X"5F",X"95",X"90",X"00",X"3F",X"99",X"99",X"00",X"5F",X"99",X"90",
		X"00",X"5F",X"99",X"99",X"00",X"59",X"99",X"99",X"00",X"59",X"99",X"99",X"00",X"55",X"99",X"99",
		X"00",X"95",X"99",X"99",X"00",X"95",X"99",X"99",X"00",X"E9",X"99",X"99",X"00",X"E9",X"93",X"99",
		X"00",X"EE",X"35",X"99",X"00",X"EE",X"55",X"99",X"00",X"AE",X"55",X"99",X"00",X"AA",X"4E",X"99",
		X"00",X"0A",X"4E",X"90",X"00",X"0A",X"AA",X"90",X"00",X"00",X"33",X"00",X"00",X"00",X"53",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"B5",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B5",X"00",X"00",X"00",X"BB",X"0F",X"00",
		X"00",X"BB",X"0F",X"00",X"00",X"B5",X"0F",X"00",X"00",X"BB",X"0F",X"00",X"00",X"55",X"00",X"00",
		X"00",X"5B",X"00",X"00",X"00",X"55",X"B0",X"00",X"00",X"55",X"B0",X"00",X"00",X"BB",X"B5",X"00",
		X"00",X"F5",X"55",X"00",X"00",X"FF",X"5B",X"00",X"0F",X"55",X"5E",X"00",X"0F",X"55",X"EB",X"00",
		X"0F",X"BB",X"BE",X"00",X"0F",X"BB",X"E5",X"00",X"0F",X"55",X"5E",X"00",X"00",X"55",X"5B",X"00",
		X"00",X"F5",X"5B",X"00",X"00",X"FF",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"B0",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"5B",X"B0",X"00",X"00",X"55",X"B0",X"00",
		X"00",X"55",X"B0",X"00",X"00",X"BF",X"B0",X"00",X"00",X"55",X"5B",X"00",X"00",X"F5",X"B5",X"00",
		X"00",X"FF",X"55",X"00",X"00",X"F5",X"B5",X"00",X"5B",X"BB",X"BB",X"00",X"5B",X"FB",X"BB",X"00",
		X"BB",X"55",X"5F",X"00",X"BB",X"B5",X"0B",X"00",X"BB",X"5B",X"0B",X"00",X"B5",X"55",X"00",X"00",
		X"F5",X"F5",X"00",X"00",X"55",X"F5",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"5F",X"00",X"00",
		X"55",X"5F",X"00",X"00",X"FB",X"5B",X"00",X"00",X"F5",X"05",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"93",X"00",
		X"90",X"99",X"99",X"00",X"99",X"AA",X"AA",X"00",X"99",X"EA",X"EA",X"09",X"99",X"F9",X"9F",X"99",
		X"99",X"5F",X"FF",X"9A",X"AA",X"99",X"99",X"95",X"57",X"99",X"FF",X"55",X"F7",X"99",X"FF",X"44",
		X"75",X"95",X"FF",X"94",X"53",X"99",X"9F",X"59",X"53",X"99",X"FF",X"59",X"53",X"99",X"FF",X"59",
		X"55",X"99",X"FF",X"59",X"55",X"95",X"FF",X"59",X"55",X"95",X"55",X"59",X"53",X"95",X"FF",X"95",
		X"73",X"3F",X"AF",X"95",X"33",X"3F",X"0A",X"55",X"35",X"3F",X"0A",X"95",X"73",X"FF",X"3A",X"94",
		X"33",X"F9",X"FF",X"4E",X"0E",X"EA",X"3A",X"EA",X"0A",X"AA",X"90",X"AA",X"5F",X"0A",X"90",X"00",
		X"99",X"0A",X"90",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",X"09",X"99",X"00",X"99",X"99",X"99",
		X"99",X"99",X"99",X"F5",X"EE",X"EE",X"EE",X"EE",X"BB",X"BB",X"BB",X"BB",X"44",X"45",X"99",X"5F",
		X"77",X"77",X"99",X"99",X"33",X"59",X"55",X"9B",X"55",X"53",X"FF",X"B5",X"5F",X"39",X"FF",X"99",
		X"FE",X"99",X"FF",X"99",X"99",X"99",X"FF",X"99",X"59",X"93",X"FF",X"99",X"59",X"93",X"FF",X"99",
		X"59",X"93",X"FF",X"99",X"59",X"93",X"FF",X"99",X"99",X"93",X"FF",X"99",X"FF",X"93",X"FF",X"99",
		X"55",X"93",X"FF",X"99",X"55",X"59",X"FF",X"55",X"33",X"59",X"55",X"95",X"77",X"77",X"99",X"99",
		X"F4",X"45",X"99",X"55",X"BF",X"BB",X"BB",X"BB",X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",
		X"E1",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"BE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",
		X"5E",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"31",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",
		X"BF",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"CC",X"99",X"99",X"90",
		X"BB",X"99",X"99",X"99",X"96",X"CC",X"CC",X"C9",X"9C",X"CA",X"BE",X"BC",X"5A",X"AE",X"AC",X"BC",
		X"AA",X"BB",X"EB",X"C9",X"9A",X"EA",X"BE",X"C5",X"EB",X"BA",X"BB",X"C9",X"BE",X"BA",X"BB",X"9C",
		X"BB",X"BA",X"BB",X"BC",X"EE",X"EA",X"BB",X"EC",X"55",X"5A",X"BB",X"BC",X"BB",X"BA",X"B5",X"EC",
		X"BB",X"BA",X"BB",X"BC",X"6F",X"BA",X"5B",X"9C",X"B6",X"BA",X"BB",X"C9",X"9B",X"BA",X"FB",X"C5",
		X"9C",X"BB",X"BB",X"C0",X"5C",X"FB",X"FF",X"BC",X"BC",X"CB",X"BB",X"BC",X"B6",X"BC",X"CC",X"C9",
		X"BB",X"99",X"99",X"90",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"01",X"79",X"00",X"99",
		X"01",X"7A",X"DD",X"99",X"09",X"77",X"9D",X"99",X"09",X"67",X"DA",X"99",X"59",X"97",X"DD",X"90",
		X"EE",X"97",X"DD",X"59",X"EE",X"97",X"DD",X"59",X"FE",X"97",X"DD",X"59",X"EE",X"27",X"DD",X"59",
		X"59",X"76",X"DD",X"50",X"09",X"67",X"DA",X"00",X"09",X"77",X"AD",X"00",X"01",X"67",X"DD",X"00",
		X"01",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"F0",X"9A",X"AA",X"AA",
		X"F5",X"7A",X"99",X"99",X"F9",X"AA",X"99",X"99",X"F9",X"EE",X"99",X"99",X"09",X"EA",X"99",X"A3",
		X"09",X"55",X"3A",X"33",X"F3",X"99",X"53",X"F9",X"39",X"93",X"7A",X"59",X"09",X"3A",X"AA",X"59",
		X"59",X"AA",X"AA",X"59",X"59",X"AF",X"99",X"59",X"59",X"FF",X"99",X"59",X"59",X"FF",X"55",X"09",
		X"59",X"FF",X"AA",X"F9",X"59",X"EF",X"AA",X"59",X"59",X"EE",X"AA",X"59",X"59",X"EE",X"AA",X"59",
		X"39",X"9E",X"EA",X"59",X"FA",X"99",X"5E",X"59",X"09",X"AE",X"EE",X"FA",X"09",X"EA",X"99",X"AA",
		X"F9",X"5E",X"99",X"EE",X"F9",X"EE",X"99",X"99",X"F5",X"AA",X"99",X"99",X"F0",X"9F",X"99",X"99",
		X"00",X"39",X"D9",X"D9",X"00",X"D0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",
		X"99",X"3A",X"99",X"00",X"99",X"99",X"99",X"F0",X"99",X"99",X"99",X"F0",X"99",X"99",X"9A",X"F0",
		X"AA",X"A7",X"99",X"F0",X"AA",X"AA",X"99",X"F0",X"AA",X"AA",X"99",X"F0",X"AA",X"94",X"9F",X"F0",
		X"AA",X"4A",X"9F",X"F0",X"AA",X"AA",X"9F",X"F0",X"AA",X"9A",X"9F",X"F0",X"AA",X"49",X"9F",X"F0",
		X"AA",X"AA",X"9F",X"F0",X"AA",X"49",X"9F",X"F0",X"AA",X"9A",X"9F",X"F0",X"AA",X"AA",X"9F",X"F0",
		X"EA",X"49",X"9F",X"F0",X"AE",X"A4",X"99",X"F0",X"EE",X"EA",X"99",X"F0",X"EE",X"EE",X"99",X"F0",
		X"99",X"99",X"9A",X"F0",X"99",X"99",X"99",X"F0",X"99",X"99",X"99",X"F0",X"D9",X"3A",X"99",X"00",
		X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"99",X"99",X"E9",
		X"99",X"EE",X"AA",X"AA",X"FF",X"AA",X"EE",X"99",X"FE",X"99",X"55",X"99",X"E9",X"99",X"99",X"99",
		X"49",X"99",X"39",X"99",X"69",X"04",X"39",X"A3",X"99",X"49",X"E9",X"EA",X"9A",X"A9",X"99",X"EE",
		X"99",X"99",X"99",X"EA",X"9A",X"49",X"99",X"AE",X"9A",X"9A",X"99",X"EA",X"9A",X"4A",X"99",X"EE",
		X"9A",X"AA",X"99",X"EA",X"9A",X"AA",X"99",X"EE",X"9E",X"49",X"99",X"E3",X"69",X"E4",X"39",X"3B",
		X"40",X"9E",X"39",X"99",X"E9",X"99",X"99",X"99",X"FE",X"99",X"55",X"99",X"FF",X"AA",X"EE",X"99",
		X"99",X"AE",X"AA",X"3A",X"09",X"99",X"99",X"A9",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",
		X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"90",X"09",X"99",X"09",X"09",X"22",X"22",X"99",X"99",X"92",X"22",
		X"99",X"99",X"92",X"22",X"21",X"33",X"92",X"22",X"13",X"A3",X"92",X"22",X"71",X"AA",X"92",X"22",
		X"13",X"FF",X"92",X"22",X"22",X"22",X"92",X"22",X"29",X"27",X"92",X"22",X"37",X"44",X"92",X"22",
		X"71",X"44",X"92",X"22",X"11",X"74",X"92",X"22",X"11",X"44",X"92",X"22",X"11",X"44",X"92",X"22",
		X"99",X"74",X"92",X"22",X"77",X"47",X"92",X"22",X"14",X"74",X"92",X"22",X"11",X"77",X"92",X"22",
		X"74",X"74",X"92",X"22",X"37",X"77",X"92",X"22",X"39",X"27",X"92",X"22",X"D3",X"22",X"92",X"22",
		X"13",X"FF",X"92",X"22",X"71",X"22",X"92",X"22",X"13",X"A2",X"92",X"22",X"21",X"33",X"92",X"22",
		X"99",X"00",X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"93",X"33",X"00",X"00",
		X"03",X"99",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",
		X"03",X"90",X"00",X"00",X"33",X"33",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"33",X"33",X"00",X"00",X"03",X"90",X"00",X"00",
		X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"99",X"00",X"00",
		X"93",X"33",X"00",X"00",X"33",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"90",X"99",
		X"90",X"09",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"DD",X"22",X"22",X"22",
		X"11",X"11",X"99",X"99",X"11",X"99",X"33",X"11",X"F7",X"99",X"11",X"19",X"11",X"99",X"7D",X"99",
		X"11",X"93",X"77",X"33",X"EE",X"93",X"77",X"33",X"97",X"93",X"77",X"33",X"97",X"93",X"77",X"33",
		X"97",X"93",X"77",X"33",X"97",X"93",X"77",X"33",X"97",X"93",X"77",X"33",X"7F",X"9F",X"77",X"33",
		X"DD",X"F3",X"75",X"33",X"EE",X"99",X"F7",X"99",X"11",X"99",X"11",X"11",X"11",X"99",X"33",X"11",
		X"77",X"77",X"99",X"99",X"5F",X"2A",X"22",X"22",X"22",X"22",X"25",X"22",X"00",X"00",X"22",X"22",
		X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"F2",X"00",X"00",X"00",
		X"F2",X"00",X"00",X"00",X"F2",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"90",X"00",X"00",X"09",X"00",X"00",X"09",X"00",X"00",X"00",X"99",X"90",X"00",X"90",
		X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"99",X"99",X"99",X"99",X"90",X"99",X"90",X"09",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",
		X"55",X"5E",X"00",X"00",X"55",X"55",X"05",X"00",X"55",X"50",X"F5",X"05",X"55",X"55",X"F5",X"55",
		X"55",X"E5",X"FF",X"55",X"55",X"5E",X"5F",X"55",X"5F",X"55",X"55",X"E5",X"F5",X"55",X"55",X"55",
		X"55",X"55",X"F5",X"55",X"55",X"5E",X"55",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"55",X"55",
		X"55",X"5F",X"F5",X"55",X"FF",X"F5",X"55",X"E5",X"55",X"F5",X"55",X"5E",X"55",X"5F",X"55",X"5E",
		X"55",X"F5",X"F5",X"55",X"55",X"5F",X"55",X"55",X"55",X"5F",X"55",X"55",X"55",X"55",X"55",X"55",
		X"55",X"55",X"55",X"55",X"5F",X"55",X"5F",X"55",X"55",X"55",X"F5",X"55",X"55",X"55",X"F5",X"55",
		X"5F",X"5F",X"FF",X"55",X"F5",X"F5",X"F5",X"55",X"55",X"5F",X"5F",X"55",X"55",X"EF",X"55",X"55",
		X"55",X"5E",X"55",X"55",X"53",X"55",X"55",X"55",X"53",X"55",X"05",X"53",X"33",X"55",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"F3",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"39",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"90",X"00",X"90",X"90",X"90",X"00",
		X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"90",
		X"90",X"90",X"90",X"90",X"90",X"90",X"90",X"00",X"90",X"90",X"90",X"00",X"00",X"90",X"90",X"00",
		X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"00",X"90",X"90",X"00",X"09",X"09",X"09",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",
		X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"00",
		X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",
		X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",
		X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",X"20",X"10",X"90",X"00",
		X"00",X"19",X"00",X"00",X"00",X"00",X"11",X"00",X"01",X"00",X"11",X"00",X"11",X"19",X"90",X"00",
		X"00",X"9D",X"00",X"00",X"00",X"9D",X"00",X"00",X"00",X"11",X"90",X"00",X"00",X"19",X"99",X"00",
		X"00",X"01",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"19",X"02",X"00",
		X"00",X"19",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"0F",X"FD",X"00",X"09",X"00",X"0F",X"00",X"99",X"0D",X"90",X"11",X"11",X"00",X"F0",X"11",
		X"11",X"0F",X"90",X"19",X"00",X"D0",X"09",X"90",X"00",X"DD",X"F0",X"00",X"01",X"1D",X"D1",X"02",
		X"01",X"11",X"01",X"00",X"00",X"11",X"01",X"00",X"00",X"00",X"09",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"22",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"19",X"00",X"00",X"00",X"11",X"10",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"90",X"00",X"60",X"00",X"11",X"0F",X"66",
		X"00",X"00",X"00",X"09",X"00",X"66",X"F0",X"00",X"44",X"00",X"00",X"FF",X"44",X"11",X"00",X"FF",
		X"41",X"11",X"66",X"00",X"99",X"66",X"00",X"66",X"00",X"10",X"66",X"0F",X"00",X"11",X"66",X"06",
		X"00",X"11",X"66",X"06",X"00",X"14",X"06",X"66",X"00",X"16",X"60",X"06",X"00",X"44",X"60",X"11",
		X"00",X"04",X"11",X"15",X"04",X"44",X"11",X"15",X"44",X"11",X"00",X"19",X"09",X"44",X"19",X"99",
		X"00",X"44",X"19",X"91",X"00",X"04",X"91",X"41",X"00",X"40",X"91",X"40",X"00",X"99",X"49",X"00",
		X"00",X"90",X"49",X"00",X"00",X"00",X"49",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"90",X"00",
		X"04",X"94",X"00",X"00",X"04",X"40",X"09",X"00",X"04",X"41",X"99",X"00",X"04",X"41",X"04",X"00",
		X"01",X"11",X"40",X"00",X"01",X"11",X"04",X"00",X"91",X"14",X"40",X"00",X"01",X"11",X"00",X"00",
		X"11",X"01",X"00",X"00",X"11",X"01",X"00",X"00",X"11",X"11",X"00",X"00",X"51",X"01",X"00",X"00",
		X"65",X"61",X"44",X"00",X"06",X"00",X"11",X"00",X"00",X"00",X"04",X"00",X"60",X"00",X"11",X"00",
		X"06",X"66",X"14",X"00",X"00",X"66",X"44",X"00",X"69",X"00",X"11",X"00",X"09",X"00",X"11",X"40",
		X"00",X"66",X"11",X"44",X"F0",X"00",X"04",X"44",X"00",X"00",X"66",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"60",X"11",X"99",X"00",X"06",X"01",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"01",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"03",X"00",X"00",X"33",X"00",X"00",
		X"00",X"33",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"43",X"00",X"00",X"00",X"43",X"00",X"39",
		X"00",X"64",X"00",X"39",X"00",X"66",X"39",X"00",X"00",X"66",X"39",X"00",X"00",X"36",X"33",X"00",
		X"00",X"16",X"61",X"00",X"00",X"6F",X"13",X"00",X"00",X"FF",X"39",X"00",X"00",X"6F",X"39",X"00",
		X"00",X"4F",X"39",X"00",X"00",X"66",X"33",X"00",X"00",X"11",X"31",X"00",X"03",X"11",X"36",X"00",
		X"00",X"31",X"13",X"00",X"03",X"31",X"13",X"00",X"00",X"11",X"11",X"00",X"00",X"31",X"33",X"00",
		X"00",X"33",X"93",X"00",X"00",X"39",X"39",X"00",X"00",X"30",X"13",X"00",X"00",X"00",X"13",X"00",
		X"00",X"09",X"00",X"00",X"00",X"99",X"00",X"90",X"00",X"61",X"00",X"99",X"00",X"91",X"09",X"00",
		X"00",X"61",X"99",X"00",X"00",X"69",X"96",X"00",X"69",X"64",X"99",X"00",X"11",X"19",X"19",X"99",
		X"31",X"99",X"99",X"99",X"09",X"99",X"99",X"99",X"93",X"11",X"99",X"99",X"63",X"66",X"99",X"99",
		X"66",X"6F",X"16",X"99",X"66",X"FF",X"13",X"90",X"16",X"6F",X"66",X"00",X"06",X"FF",X"31",X"00",
		X"01",X"FF",X"F6",X"00",X"00",X"FF",X"69",X"00",X"66",X"4F",X"19",X"90",X"06",X"FF",X"66",X"90",
		X"33",X"F6",X"99",X"00",X"06",X"66",X"11",X"00",X"66",X"1F",X"16",X"00",X"66",X"66",X"36",X"00",
		X"19",X"66",X"66",X"90",X"99",X"99",X"69",X"90",X"09",X"99",X"99",X"99",X"03",X"99",X"99",X"90",
		X"06",X"10",X"09",X"00",X"66",X"90",X"90",X"09",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"09",X"90",X"00",X"99",X"99",X"00",
		X"00",X"19",X"96",X"00",X"00",X"99",X"66",X"00",X"99",X"49",X"11",X"00",X"19",X"99",X"33",X"39",
		X"10",X"99",X"39",X"33",X"90",X"91",X"99",X"93",X"39",X"11",X"31",X"66",X"33",X"66",X"91",X"61",
		X"33",X"36",X"99",X"19",X"33",X"66",X"11",X"99",X"00",X"31",X"63",X"90",X"00",X"64",X"16",X"90",
		X"00",X"66",X"99",X"03",X"00",X"36",X"99",X"33",X"00",X"66",X"33",X"30",X"00",X"36",X"91",X"00",
		X"30",X"34",X"93",X"00",X"03",X"64",X"93",X"03",X"63",X"69",X"99",X"33",X"69",X"33",X"91",X"33",
		X"99",X"99",X"66",X"30",X"00",X"93",X"16",X"90",X"91",X"96",X"11",X"99",X"03",X"99",X"99",X"99",
		X"03",X"09",X"99",X"99",X"06",X"00",X"03",X"99",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",
		X"00",X"99",X"99",X"00",X"00",X"93",X"99",X"00",X"04",X"93",X"33",X"00",X"19",X"33",X"93",X"00",
		X"00",X"93",X"33",X"00",X"00",X"19",X"99",X"00",X"01",X"93",X"36",X"90",X"03",X"66",X"66",X"90",
		X"03",X"19",X"91",X"39",X"06",X"31",X"99",X"99",X"33",X"96",X"99",X"90",X"09",X"31",X"39",X"00",
		X"00",X"99",X"39",X"00",X"30",X"33",X"33",X"00",X"99",X"66",X"93",X"00",X"33",X"99",X"33",X"00",
		X"93",X"19",X"33",X"00",X"39",X"19",X"39",X"00",X"33",X"99",X"33",X"00",X"93",X"93",X"33",X"00",
		X"99",X"93",X"93",X"30",X"99",X"93",X"39",X"39",X"99",X"93",X"99",X"33",X"90",X"99",X"93",X"99",
		X"00",X"39",X"39",X"99",X"00",X"90",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"09",X"33",X"00",X"00",X"99",X"33",X"00",X"00",X"03",X"33",X"00",
		X"00",X"33",X"30",X"00",X"00",X"33",X"90",X"00",X"00",X"33",X"90",X"00",X"00",X"99",X"33",X"99",
		X"00",X"33",X"33",X"33",X"00",X"33",X"33",X"00",X"00",X"33",X"33",X"00",X"03",X"33",X"93",X"03",
		X"33",X"39",X"93",X"00",X"33",X"33",X"33",X"00",X"03",X"33",X"33",X"00",X"00",X"33",X"33",X"00",
		X"00",X"93",X"33",X"00",X"00",X"33",X"93",X"00",X"00",X"33",X"99",X"00",X"00",X"33",X"09",X"00",
		X"00",X"03",X"30",X"30",X"00",X"03",X"33",X"30",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"09",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"09",X"00",X"00",X"30",X"39",X"00",X"30",X"50",X"33",X"00",X"30",X"50",X"33",X"00",
		X"00",X"55",X"30",X"00",X"00",X"35",X"53",X"00",X"03",X"3F",X"F5",X"33",X"33",X"33",X"F3",X"30",
		X"55",X"99",X"93",X"90",X"00",X"99",X"F3",X"00",X"33",X"39",X"F3",X"00",X"03",X"99",X"3F",X"00",
		X"09",X"39",X"3F",X"09",X"00",X"99",X"35",X"30",X"00",X"99",X"F5",X"00",X"03",X"33",X"33",X"00",
		X"59",X"53",X"F3",X"30",X"33",X"33",X"33",X"03",X"00",X"55",X"30",X"00",X"00",X"50",X"03",X"00",
		X"00",X"50",X"33",X"00",X"00",X"00",X"30",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"90",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"FF",X"44",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"FF",X"66",X"00",
		X"00",X"FF",X"16",X"00",X"00",X"F5",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"FF",X"44",X"00",
		X"00",X"FF",X"66",X"00",X"00",X"55",X"46",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"07",X"55",X"11",X"00",X"77",X"FF",X"66",X"00",
		X"77",X"FF",X"11",X"01",X"07",X"55",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"75",X"55",X"00",X"00",X"77",X"FF",X"11",X"00",X"77",X"FF",X"66",X"00",
		X"77",X"FF",X"11",X"01",X"75",X"55",X"61",X"02",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"75",X"55",X"00",X"00",X"77",X"FF",X"66",X"40",X"77",X"FF",X"44",X"00",
		X"77",X"FF",X"64",X"06",X"75",X"55",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"49",X"69",X"00",X"00",X"04",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"40",X"00",X"00",X"00",X"69",X"00",X"00",X"00",X"46",X"04",X"00",X"00",X"04",X"90",X"00",
		X"00",X"04",X"90",X"00",X"00",X"09",X"90",X"00",X"00",X"69",X"40",X"00",X"00",X"09",X"40",X"00",
		X"00",X"09",X"04",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"33",X"0F",X"00",X"00",X"05",X"FF",X"00",
		X"00",X"4F",X"35",X"00",X"00",X"44",X"43",X"00",X"00",X"44",X"FF",X"00",X"00",X"F4",X"55",X"00",
		X"00",X"44",X"3F",X"00",X"00",X"66",X"44",X"00",X"00",X"46",X"44",X"00",X"00",X"54",X"54",X"00",
		X"00",X"54",X"00",X"00",X"00",X"FF",X"05",X"00",X"00",X"FF",X"45",X"00",X"00",X"05",X"4F",X"00",
		X"00",X"05",X"F4",X"00",X"00",X"04",X"00",X"00",X"00",X"F4",X"00",X"00",X"00",X"54",X"00",X"00",
		X"00",X"04",X"06",X"00",X"00",X"0F",X"00",X"00",X"00",X"4F",X"00",X"00",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"E5",X"50",X"00",X"00",X"33",X"5F",X"00",X"00",X"F5",X"FF",X"00",
		X"00",X"4F",X"35",X"00",X"00",X"45",X"43",X"00",X"00",X"44",X"FF",X"00",X"00",X"F4",X"55",X"00",
		X"00",X"FF",X"3F",X"00",X"00",X"FF",X"53",X"00",X"00",X"FF",X"F4",X"00",X"00",X"5F",X"54",X"00",
		X"00",X"54",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"FF",X"45",X"00",X"00",X"F5",X"4F",X"00",
		X"00",X"F5",X"F4",X"00",X"00",X"F3",X"F3",X"00",X"00",X"FE",X"00",X"00",X"00",X"5F",X"F0",X"00",
		X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"50",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"35",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"E5",X"5F",X"00",X"00",X"33",X"5F",X"00",X"00",X"F5",X"55",X"00",
		X"03",X"FF",X"35",X"00",X"00",X"55",X"53",X"00",X"05",X"55",X"5F",X"00",X"55",X"55",X"55",X"00",
		X"55",X"53",X"3F",X"00",X"05",X"55",X"53",X"00",X"00",X"5F",X"5F",X"00",X"00",X"5F",X"53",X"00",
		X"00",X"55",X"55",X"00",X"00",X"55",X"F5",X"00",X"00",X"FF",X"F5",X"00",X"00",X"F5",X"FF",X"00",
		X"00",X"F5",X"FF",X"00",X"00",X"F3",X"F3",X"00",X"00",X"FE",X"EE",X"00",X"00",X"5F",X"F5",X"00",
		X"00",X"55",X"55",X"00",X"00",X"FF",X"55",X"00",X"00",X"5F",X"5F",X"00",X"00",X"FF",X"50",X"00",
		X"00",X"55",X"00",X"53",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"EE",X"E0",X"00",X"00",X"55",X"55",X"00",
		X"00",X"5F",X"F5",X"00",X"00",X"5F",X"3F",X"00",X"00",X"5F",X"F5",X"00",X"00",X"3E",X"F5",X"00",
		X"EE",X"EF",X"55",X"00",X"E5",X"5F",X"55",X"00",X"E5",X"FF",X"55",X"00",X"55",X"5F",X"F5",X"00",
		X"50",X"5F",X"F3",X"00",X"5F",X"FF",X"5F",X"00",X"55",X"5F",X"5F",X"00",X"55",X"5F",X"5F",X"00",
		X"55",X"FF",X"5F",X"00",X"E5",X"FF",X"FF",X"00",X"E5",X"FF",X"F3",X"00",X"E3",X"F5",X"FF",X"00",
		X"33",X"F3",X"55",X"00",X"00",X"53",X"55",X"00",X"00",X"35",X"FF",X"00",X"30",X"55",X"F5",X"30",
		X"30",X"55",X"F5",X"00",X"00",X"55",X"55",X"33",X"00",X"55",X"EE",X"53",X"00",X"FE",X"00",X"F3",
		X"00",X"33",X"00",X"F5",X"00",X"E0",X"30",X"55",X"00",X"00",X"03",X"50",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"1A",X"00",X"00",X"00",X"66",X"64",X"00",X"00",X"04",X"06",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"0A",X"11",X"06",X"00",
		X"0A",X"66",X"00",X"00",X"44",X"44",X"00",X"00",X"64",X"00",X"00",X"00",X"66",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"16",X"64",X"04",X"00",X"0A",X"06",X"00",X"00",X"A6",X"00",X"00",X"00",
		X"61",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"11",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"26",X"66",X"00",X"00",X"00",X"44",X"00",X"00",
		X"00",X"61",X"00",X"00",X"00",X"16",X"00",X"00",X"02",X"01",X"00",X"00",X"66",X"00",X"60",X"00",
		X"44",X"10",X"06",X"00",X"02",X"06",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"44",X"66",X"00",X"00",X"66",X"41",X"04",X"00",X"44",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"0A",X"60",X"00",X"00",X"06",X"06",X"06",X"00",X"04",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"04",X"00",X"00",X"00",
		X"44",X"00",X"00",X"00",X"66",X"41",X"04",X"00",X"44",X"66",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"02",X"06",X"00",X"06",X"44",X"10",X"00",X"60",
		X"66",X"00",X"60",X"00",X"02",X"01",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"00",X"00",X"00",X"26",X"66",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"06",X"00",
		X"00",X"11",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"61",X"00",X"00",X"00",
		X"A6",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"16",X"61",X"04",X"00",X"44",X"06",X"00",X"00",
		X"66",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"44",X"44",X"00",X"00",X"0A",X"00",X"00",X"00",
		X"0A",X"11",X"06",X"00",X"06",X"66",X"00",X"00",X"66",X"44",X"60",X"00",X"44",X"00",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"04",X"06",X"00",X"00",X"66",X"64",X"00",X"00",X"1A",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"03",
		X"99",X"79",X"00",X"00",X"96",X"79",X"00",X"00",X"06",X"77",X"90",X"00",X"04",X"77",X"99",X"00",
		X"09",X"17",X"99",X"00",X"09",X"12",X"99",X"00",X"09",X"12",X"99",X"00",X"D9",X"22",X"D9",X"00",
		X"11",X"27",X"DD",X"00",X"11",X"77",X"DD",X"00",X"57",X"DD",X"AD",X"00",X"90",X"77",X"0A",X"00",
		X"90",X"77",X"90",X"00",X"00",X"D7",X"EE",X"00",X"00",X"DD",X"EE",X"00",X"00",X"00",X"EE",X"00",
		X"00",X"00",X"EE",X"00",X"00",X"00",X"E5",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"90",
		X"00",X"00",X"00",X"90",X"00",X"00",X"A0",X"90",X"00",X"00",X"A0",X"90",X"00",X"00",X"DA",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"D2",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0D",X"09",
		X"00",X"00",X"0D",X"F9",X"00",X"00",X"DD",X"99",X"00",X"00",X"DD",X"99",X"00",X"00",X"DA",X"99",
		X"00",X"00",X"AE",X"00",X"00",X"00",X"AE",X"90",X"00",X"00",X"DA",X"09",X"00",X"70",X"DD",X"90",
		X"00",X"77",X"AD",X"90",X"00",X"67",X"AD",X"09",X"00",X"06",X"AD",X"20",X"00",X"07",X"DD",X"29",
		X"00",X"07",X"DD",X"20",X"00",X"02",X"97",X"00",X"00",X"11",X"99",X"00",X"00",X"15",X"09",X"00",
		X"00",X"1F",X"90",X"00",X"00",X"11",X"09",X"00",X"00",X"11",X"90",X"00",X"00",X"90",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"09",X"97",X"00",X"00",X"09",X"11",X"00",X"00",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"00",X"F0",X"60",X"0B",X"06",X"00",X"60",
		X"BB",X"66",X"66",X"00",X"00",X"64",X"A4",X"AA",X"00",X"64",X"44",X"EE",X"4B",X"55",X"AF",X"0B",
		X"EF",X"55",X"AF",X"00",X"BF",X"56",X"99",X"EE",X"B0",X"15",X"B0",X"EE",X"44",X"F1",X"00",X"EB",
		X"00",X"FF",X"50",X"1E",X"0F",X"FF",X"FF",X"0E",X"44",X"FF",X"F0",X"55",X"01",X"FF",X"11",X"F5",
		X"44",X"FF",X"F0",X"55",X"06",X"FF",X"11",X"55",X"00",X"FF",X"FF",X"5B",X"F4",X"11",X"00",X"EE",
		X"44",X"91",X"00",X"BE",X"44",X"69",X"99",X"EE",X"E0",X"66",X"0A",X"BE",X"00",X"00",X"01",X"EB",
		X"00",X"00",X"01",X"EE",X"00",X"B0",X"00",X"AF",X"B0",X"99",X"69",X"00",X"BB",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"90",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"AA",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"A1",
		X"00",X"00",X"00",X"11",X"00",X"06",X"00",X"1A",X"00",X"00",X"10",X"1A",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"96",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"60",X"66",X"00",X"00",X"66",X"64",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"4E",
		X"00",X"00",X"00",X"11",X"00",X"00",X"F0",X"51",X"00",X"00",X"FF",X"61",X"00",X"60",X"0F",X"51",
		X"00",X"00",X"4F",X"11",X"00",X"01",X"64",X"F5",X"00",X"00",X"6F",X"F1",X"00",X"00",X"41",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"11",X"60",X"00",X"00",
		X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"64",X"00",X"00",X"00",X"61",X"00",X"10",X"00",
		X"16",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"11",X"00",X"00",X"66",X"10",X"00",X"B0",
		X"66",X"00",X"00",X"00",X"61",X"0B",X"BB",X"00",X"FF",X"BB",X"BE",X"00",X"11",X"BB",X"11",X"00",
		X"00",X"60",X"11",X"FF",X"00",X"00",X"44",X"FF",X"00",X"00",X"66",X"FF",X"00",X"11",X"06",X"FF",
		X"00",X"10",X"00",X"1F",X"00",X"00",X"66",X"11",X"00",X"00",X"66",X"91",X"00",X"00",X"66",X"66",
		X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"11",X"00",X"01",X"00",X"11",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"01",X"00",X"00",X"0B",X"01",X"00",
		X"00",X"0B",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AB",X"00",X"00",X"00",X"AB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"61",X"44",X"00",X"00",X"66",X"11",X"60",X"00",X"66",X"66",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"16",X"11",X"11",X"BE",X"66",X"00",X"00",X"00",X"61",X"11",X"00",X"00",X"66",X"10",X"00",X"00",
		X"11",X"66",X"00",X"00",X"11",X"00",X"00",X"00",X"01",X"10",X"00",X"00",X"91",X"11",X"00",X"00",
		X"06",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"06",X"00",X"00",X"60",X"00",X"00",X"00",
		X"66",X"00",X"10",X"00",X"06",X"00",X"00",X"00",X"06",X"10",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"B0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"66",
		X"00",X"01",X"00",X"61",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",
		X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"91",X"00",X"00",X"66",X"11",X"00",X"10",X"00",X"1F",
		X"06",X"11",X"06",X"FF",X"00",X"00",X"66",X"FF",X"00",X"00",X"44",X"FF",X"00",X"60",X"11",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"06",X"10",X"10",X"00",X"06",X"00",X"00",X"00",X"66",X"00",X"10",X"00",
		X"60",X"00",X"00",X"00",X"60",X"06",X"00",X"00",X"60",X"00",X"00",X"00",X"06",X"00",X"00",X"00",
		X"91",X"11",X"00",X"00",X"01",X"10",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"66",X"00",X"00",
		X"66",X"10",X"00",X"00",X"61",X"11",X"00",X"00",X"66",X"00",X"00",X"00",X"16",X"11",X"11",X"BE",
		X"FF",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"11",X"60",X"00",X"61",X"44",X"00",X"00",
		X"00",X"00",X"41",X"6F",X"00",X"00",X"6F",X"61",X"00",X"01",X"64",X"66",X"00",X"00",X"4F",X"16",
		X"00",X"60",X"0F",X"66",X"00",X"00",X"FF",X"66",X"00",X"00",X"F0",X"55",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"4E",X"00",X"00",X"00",X"44",X"00",X"00",X"66",X"64",X"00",X"00",X"60",X"66",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"01",X"96",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"1A",X"00",X"06",X"00",X"1A",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"A1",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"60",X"00",X"10",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"BB",X"11",X"00",X"FF",X"BB",X"BE",X"00",X"61",X"0B",X"00",X"00",X"66",X"00",X"00",X"00",
		X"61",X"16",X"00",X"00",X"66",X"11",X"00",X"00",X"66",X"00",X"00",X"00",X"16",X"00",X"60",X"00",
		X"61",X"00",X"16",X"00",X"64",X"11",X"00",X"00",X"66",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"60",X"00",X"00",X"19",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"96",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",
		X"00",X"00",X"00",X"06",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"00",X"03",
		X"00",X"00",X"00",X"33",X"00",X"00",X"F0",X"53",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"03",
		X"00",X"00",X"4F",X"13",X"00",X"00",X"64",X"03",X"00",X"00",X"60",X"03",X"00",X"00",X"41",X"33",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"61",X"00",X"00",X"00",X"19",X"00",X"00",X"00",X"11",X"60",X"00",X"00",
		X"11",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"64",X"11",X"00",X"00",X"63",X"00",X"16",X"00",
		X"33",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"33",X"11",X"00",X"00",X"00",X"16",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"11",X"33",X"00",X"00",X"44",X"33",X"00",X"00",X"66",X"00",X"00",X"01",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"30",X"00",X"00",X"60",X"33",X"00",X"00",X"60",X"33",
		X"00",X"00",X"00",X"36",X"00",X"00",X"00",X"33",X"00",X"00",X"00",X"61",X"00",X"01",X"00",X"61",
		X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"11",X"60",X"00",X"00",X"66",X"30",X"00",X"00",X"00",X"00",X"00",
		X"00",X"01",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",
		X"33",X"33",X"00",X"00",X"33",X"03",X"00",X"00",X"31",X"10",X"00",X"00",X"31",X"01",X"00",X"00",
		X"36",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"60",X"06",X"00",X"00",X"60",X"00",X"00",X"00",
		X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"0B",X"0B",X"00",X"00",X"00",X"A0",X"00",X"0E",X"EE",X"AA",X"0A",X"45",X"99",X"00",
		X"BB",X"77",X"99",X"FB",X"A0",X"59",X"FF",X"93",X"A5",X"53",X"FF",X"F5",X"5F",X"39",X"FF",X"99",
		X"F5",X"99",X"FF",X"95",X"55",X"99",X"FF",X"F9",X"55",X"93",X"FF",X"F9",X"33",X"93",X"FF",X"F9",
		X"33",X"93",X"FF",X"F9",X"55",X"93",X"FF",X"F9",X"55",X"93",X"FF",X"F9",X"F5",X"93",X"FF",X"95",
		X"5F",X"93",X"FF",X"99",X"05",X"59",X"FF",X"F5",X"0B",X"59",X"FF",X"9B",X"00",X"77",X"99",X"F9",
		X"00",X"45",X"99",X"00",X"B0",X"00",X"EE",X"0A",X"0B",X"00",X"AB",X"00",X"0A",X"A0",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A0",X"00",X"A0",X"00",X"00",X"0A",X"0A",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"59",X"FF",X"A0",X"00",X"53",X"FF",X"0A",X"0A",X"39",X"FF",X"0A",
		X"A5",X"99",X"FF",X"00",X"05",X"99",X"FF",X"00",X"05",X"93",X"FF",X"00",X"03",X"93",X"FF",X"00",
		X"03",X"93",X"FF",X"00",X"05",X"93",X"FF",X"00",X"00",X"93",X"FF",X"00",X"A0",X"93",X"FF",X"0B",
		X"BA",X"93",X"FF",X"0B",X"B0",X"59",X"FF",X"0B",X"0B",X"59",X"FF",X"BB",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0B",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",
		X"00",X"AA",X"B0",X"0B",X"00",X"00",X"BB",X"00",X"0A",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",
		X"AB",X"55",X"F0",X"00",X"0B",X"99",X"FF",X"00",X"00",X"93",X"FF",X"00",X"00",X"93",X"FF",X"00",
		X"00",X"93",X"FF",X"00",X"00",X"93",X"FF",X"00",X"0B",X"93",X"FF",X"00",X"AB",X"93",X"FF",X"00",
		X"A0",X"03",X"FF",X"00",X"0A",X"00",X"FF",X"00",X"00",X"00",X"F0",X"0B",X"00",X"A0",X"00",X"0B",
		X"00",X"0A",X"00",X"0B",X"00",X"00",X"B0",X"B0",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"AA",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"0A",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"30",X"09",X"00",X"00",X"33",X"93",X"00",X"00",X"03",X"33",X"00",X"00",X"03",X"30",X"00",
		X"00",X"03",X"90",X"00",X"00",X"01",X"90",X"00",X"00",X"16",X"90",X"00",X"00",X"66",X"90",X"00",
		X"00",X"66",X"90",X"00",X"00",X"66",X"90",X"00",X"00",X"16",X"90",X"00",X"00",X"01",X"90",X"00",
		X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",
		X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",X"00",X"03",X"90",X"00",
		X"00",X"03",X"39",X"00",X"00",X"03",X"33",X"00",X"00",X"33",X"03",X"00",X"00",X"30",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",
		X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"88",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"B0",X"BB",
		X"00",X"00",X"B0",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"BB",X"00",X"00",X"BB",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",
		X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"0B",X"BB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",
		X"00",X"0B",X"B0",X"00",X"00",X"0B",X"00",X"00",X"0B",X"0B",X"00",X"00",X"0B",X"0B",X"00",X"00",
		X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",
		X"BB",X"0B",X"00",X"B0",X"BB",X"BB",X"00",X"B0",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"B0",X"00",
		X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"00",X"B0",
		X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"00",X"B0",X"BB",X"BB",X"00",X"B0",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"BB",X"BB",
		X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"00",X"00",X"BB",X"BB",X"00",X"00",X"B0",X"BB",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"0B",X"BB",X"00",X"00",X"B0",X"BB",
		X"00",X"00",X"B0",X"BB",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"B0",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"00",X"B0",X"BB",X"BB",X"00",X"B0",X"BB",X"BB",X"BB",X"B0",
		X"BB",X"BB",X"00",X"B0",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"B0",X"00",
		X"BB",X"BB",X"B0",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"B0",X"BB",X"0B",X"00",X"B0",
		X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"0B",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"B0",X"00",X"00",X"BB",X"B0",X"00",X"00",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",
		X"0B",X"0B",X"00",X"00",X"0B",X"0B",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"0B",X"B0",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"92",X"22",X"22",
		X"22",X"92",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"29",X"22",X"22",X"99",X"29",X"22",
		X"22",X"99",X"29",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",
		X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"99",X"22",X"22",
		X"22",X"A9",X"2A",X"22",X"22",X"AA",X"AA",X"22",X"22",X"AA",X"AA",X"22",X"22",X"9A",X"A9",X"22",
		X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"92",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"92",X"22",
		X"22",X"22",X"92",X"22",X"22",X"99",X"99",X"22",X"22",X"99",X"99",X"22",X"22",X"99",X"E9",X"22",
		X"22",X"99",X"E9",X"22",X"22",X"99",X"E9",X"22",X"22",X"99",X"99",X"22",X"22",X"99",X"E9",X"22",
		X"22",X"99",X"E9",X"22",X"22",X"99",X"E9",X"22",X"22",X"99",X"99",X"22",X"22",X"99",X"E9",X"22",
		X"22",X"99",X"E9",X"22",X"22",X"99",X"EE",X"22",X"22",X"99",X"99",X"22",X"22",X"22",X"92",X"22",
		X"22",X"22",X"92",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"99",X"99",X"99",X"99",X"22",X"22",X"22",X"99",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"22",X"29",X"29",X"29",X"22",
		X"22",X"92",X"92",X"22",X"29",X"29",X"29",X"22",X"22",X"92",X"92",X"22",X"29",X"9F",X"29",X"22",
		X"22",X"9F",X"92",X"22",X"29",X"EE",X"99",X"22",X"22",X"55",X"92",X"22",X"29",X"55",X"99",X"22",
		X"22",X"FF",X"92",X"22",X"29",X"5F",X"99",X"22",X"22",X"FF",X"92",X"22",X"29",X"FF",X"29",X"22",
		X"22",X"9F",X"92",X"22",X"29",X"29",X"29",X"22",X"22",X"92",X"92",X"22",X"29",X"29",X"29",X"22",
		X"22",X"92",X"92",X"22",X"99",X"99",X"99",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",
		X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",
		X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",
		X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",
		X"09",X"09",X"09",X"00",X"90",X"90",X"90",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",X"09",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"09",X"09",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"E5",X"55",X"00",X"00",X"FF",X"FF",
		X"00",X"99",X"FF",X"FF",X"00",X"FF",X"EE",X"EE",X"00",X"FF",X"99",X"99",X"00",X"FF",X"99",X"9E",
		X"00",X"F5",X"EE",X"55",X"99",X"F5",X"F5",X"99",X"00",X"F5",X"FF",X"EE",X"0F",X"55",X"FF",X"99",
		X"FF",X"53",X"EE",X"24",X"FF",X"53",X"FE",X"42",X"FF",X"53",X"FE",X"24",X"FF",X"53",X"F5",X"42",
		X"FF",X"53",X"F5",X"24",X"FF",X"53",X"FE",X"42",X"FF",X"53",X"F5",X"24",X"FF",X"53",X"FF",X"22",
		X"0F",X"55",X"FF",X"99",X"00",X"F5",X"FF",X"FF",X"99",X"F5",X"FF",X"99",X"00",X"F5",X"55",X"FF",
		X"00",X"FF",X"33",X"35",X"00",X"FF",X"33",X"33",X"00",X"FF",X"55",X"55",X"00",X"5F",X"FF",X"FF",
		X"00",X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"E9",X"99",X"99",X"00",X"55",X"55",X"55",X"00",
		X"FF",X"FF",X"FE",X"00",X"EE",X"FF",X"FE",X"00",X"EF",X"22",X"FE",X"00",X"F2",X"44",X"FE",X"00",
		X"24",X"44",X"FE",X"00",X"24",X"44",X"FE",X"00",X"24",X"44",X"FE",X"00",X"24",X"44",X"FE",X"00",
		X"24",X"44",X"FE",X"00",X"24",X"44",X"FE",X"00",X"44",X"44",X"FE",X"00",X"44",X"44",X"FE",X"00",
		X"24",X"44",X"FE",X"00",X"24",X"44",X"FE",X"00",X"24",X"44",X"FE",X"00",X"24",X"44",X"FE",X"00",
		X"24",X"44",X"FE",X"00",X"44",X"44",X"FE",X"00",X"24",X"24",X"FE",X"00",X"22",X"22",X"FE",X"00",
		X"32",X"22",X"FE",X"00",X"53",X"FF",X"FE",X"00",X"55",X"FF",X"FE",X"00",X"FF",X"FF",X"FF",X"00",
		X"FF",X"55",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"9E",X"00",
		X"00",X"99",X"99",X"0E",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"EE",
		X"00",X"94",X"55",X"EE",X"09",X"49",X"55",X"EE",X"99",X"99",X"55",X"EE",X"99",X"99",X"55",X"EE",
		X"99",X"99",X"53",X"EE",X"94",X"99",X"59",X"EE",X"49",X"99",X"99",X"EE",X"AA",X"AA",X"A9",X"99",
		X"4A",X"AA",X"F9",X"EE",X"A4",X"AA",X"F9",X"EE",X"AA",X"AA",X"F9",X"EE",X"9A",X"AA",X"FF",X"EE",
		X"99",X"AA",X"FF",X"EE",X"09",X"4A",X"FF",X"EE",X"00",X"A4",X"FF",X"EE",X"00",X"AA",X"AA",X"5E",
		X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"99",X"0E",X"00",X"00",X"9E",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"5E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"0A",X"AA",X"00",X"00",X"00",X"1A",X"00",X"00",X"99",X"11",X"00",X"00",X"00",X"11",X"00",
		X"00",X"09",X"11",X"00",X"00",X"90",X"1A",X"00",X"06",X"00",X"10",X"00",X"00",X"99",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"A0",X"00",X"00",X"00",X"10",X"00",X"00",X"90",X"1A",X"00",X"00",X"09",X"11",X"00",
		X"00",X"00",X"11",X"00",X"00",X"99",X"11",X"00",X"00",X"00",X"1A",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0E",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"99",X"00",
		X"00",X"05",X"E9",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"05",X"99",X"00",
		X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"05",X"99",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"50",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"F0",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"99",X"99",X"00",X"CC",X"99",X"99",X"90",
		X"BB",X"99",X"99",X"99",X"96",X"CC",X"CC",X"C9",X"9C",X"CA",X"BE",X"BC",X"5A",X"AE",X"AC",X"B1",
		X"AA",X"BB",X"EB",X"C9",X"9A",X"EA",X"BE",X"C1",X"EB",X"BA",X"BB",X"C9",X"BE",X"BA",X"BB",X"91",
		X"BB",X"BA",X"BB",X"BC",X"EE",X"EA",X"BB",X"EC",X"55",X"5A",X"BB",X"BC",X"BB",X"BA",X"B5",X"EC",
		X"BB",X"BA",X"BB",X"BC",X"6F",X"BA",X"5B",X"91",X"B6",X"BA",X"BB",X"C9",X"9B",X"BA",X"FB",X"C1",
		X"9C",X"BB",X"BB",X"C0",X"5C",X"FB",X"FF",X"B1",X"BC",X"CB",X"BB",X"BC",X"B6",X"BC",X"CC",X"C9",
		X"BB",X"99",X"99",X"90",X"CC",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"01",X"79",X"00",X"99",
		X"01",X"7A",X"DD",X"19",X"09",X"77",X"9D",X"91",X"09",X"67",X"DA",X"69",X"59",X"97",X"DD",X"61",
		X"EE",X"97",X"DD",X"19",X"EE",X"97",X"DD",X"59",X"FE",X"97",X"DD",X"59",X"EE",X"27",X"DD",X"19",
		X"59",X"76",X"DD",X"61",X"09",X"67",X"DA",X"60",X"09",X"77",X"AD",X"01",X"01",X"67",X"DD",X"10",
		X"01",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"99",X"00",
		X"99",X"3A",X"99",X"10",X"99",X"99",X"99",X"F0",X"99",X"99",X"99",X"10",X"99",X"99",X"9A",X"F0",
		X"AA",X"A7",X"99",X"10",X"AA",X"AA",X"99",X"F0",X"AA",X"AA",X"99",X"10",X"AA",X"94",X"9F",X"F0",
		X"AA",X"4A",X"9F",X"F0",X"AA",X"AA",X"9F",X"F0",X"AA",X"9A",X"9F",X"F0",X"AA",X"49",X"9F",X"F0",
		X"AA",X"AA",X"9F",X"F0",X"AA",X"49",X"9F",X"F0",X"AA",X"9A",X"9F",X"F0",X"AA",X"AA",X"9F",X"F0",
		X"EA",X"49",X"9F",X"F0",X"AE",X"A4",X"99",X"10",X"EE",X"EA",X"99",X"F0",X"EE",X"EE",X"99",X"10",
		X"99",X"99",X"9A",X"F0",X"99",X"99",X"99",X"10",X"99",X"99",X"99",X"F0",X"D9",X"3A",X"99",X"10",
		X"00",X"99",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EA",X"00",X"00",X"00",
		X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"33",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"16",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"61",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"67",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"09",X"00",X"90",X"99",X"99",X"00",X"99",X"99",X"99",X"99",X"99",X"99",X"99",
		X"59",X"99",X"99",X"99",X"59",X"AE",X"99",X"EE",X"59",X"EA",X"99",X"E5",X"59",X"AE",X"AE",X"99",
		X"59",X"EA",X"9A",X"9A",X"53",X"A9",X"AF",X"FF",X"39",X"99",X"9A",X"9A",X"99",X"A7",X"99",X"99",
		X"99",X"AA",X"7A",X"7A",X"FF",X"AA",X"AE",X"AE",X"99",X"A9",X"EA",X"EA",X"99",X"99",X"EE",X"AE",
		X"FF",X"9F",X"EA",X"EA",X"99",X"9F",X"EE",X"AE",X"99",X"99",X"EE",X"EA",X"FF",X"9F",X"5E",X"AE",
		X"99",X"9F",X"E5",X"EE",X"99",X"E9",X"5E",X"EE",X"FF",X"E9",X"E5",X"E5",X"99",X"EE",X"65",X"55",
		X"99",X"5E",X"AA",X"AA",X"39",X"99",X"DD",X"DD",X"53",X"AA",X"DF",X"FF",X"50",X"EE",X"DD",X"DD",
		X"50",X"5E",X"AA",X"AA",X"50",X"EE",X"EE",X"E5",X"50",X"EA",X"09",X"EE",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"DA",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"11",X"11",X"FF",X"FF",X"11",X"11",X"55",X"5F",X"11",X"11",X"BB",X"5F",X"11",X"11",X"AB",X"5F",
		X"11",X"11",X"AB",X"5F",X"11",X"19",X"AB",X"5F",X"11",X"11",X"AB",X"5F",X"22",X"22",X"AA",X"A5",
		X"91",X"22",X"99",X"95",X"29",X"22",X"99",X"95",X"09",X"22",X"FF",X"FF",X"09",X"22",X"AB",X"B5",
		X"09",X"99",X"9A",X"B5",X"01",X"11",X"9A",X"B5",X"09",X"11",X"9A",X"B5",X"02",X"22",X"9A",X"BB",
		X"09",X"11",X"9A",X"AA",X"00",X"11",X"99",X"99",X"00",X"11",X"99",X"99",X"00",X"11",X"FF",X"FF",
		X"00",X"11",X"55",X"55",X"00",X"11",X"99",X"91",X"00",X"22",X"12",X"22",X"00",X"11",X"21",X"12",
		X"00",X"11",X"11",X"11",X"00",X"11",X"11",X"22",X"00",X"11",X"11",X"22",X"00",X"11",X"19",X"99",
		X"00",X"19",X"91",X"99",X"00",X"00",X"00",X"00",X"00",X"EE",X"EE",X"99",X"00",X"99",X"99",X"90",
		X"29",X"22",X"22",X"92",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"99",X"99",X"99",X"99",
		X"22",X"22",X"22",X"92",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"33",X"33",X"23",X"33",X"99",X"92",X"99",X"99",
		X"33",X"33",X"33",X"33",X"33",X"33",X"33",X"31",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"11",X"11",X"11",X"11",X"22",X"11",X"22",X"21",X"22",X"11",X"11",X"11",X"22",X"22",
		X"11",X"11",X"99",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"11",X"11",X"91",X"11",X"11",X"11",X"92",X"29",X"12",X"11",X"99",X"99",X"21",X"22",X"99",X"99",
		X"00",X"99",X"99",X"93",X"00",X"E3",X"EE",X"99",X"00",X"33",X"33",X"33",X"00",X"19",X"91",X"99",
		X"00",X"22",X"19",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",
		X"00",X"22",X"29",X"22",X"00",X"99",X"99",X"29",X"00",X"11",X"99",X"22",X"00",X"22",X"99",X"22",
		X"00",X"22",X"99",X"22",X"00",X"22",X"33",X"22",X"00",X"22",X"EE",X"22",X"09",X"99",X"FE",X"19",
		X"02",X"12",X"FE",X"92",X"09",X"22",X"EE",X"22",X"02",X"22",X"5E",X"22",X"09",X"22",X"55",X"22",
		X"29",X"99",X"22",X"29",X"02",X"22",X"92",X"22",X"22",X"22",X"22",X"22",X"92",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"29",X"22",X"22",X"99",X"22",X"92",X"99",X"22",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",
		X"11",X"19",X"00",X"00",X"11",X"19",X"90",X"00",X"11",X"19",X"09",X"00",X"11",X"19",X"90",X"00",
		X"11",X"12",X"00",X"00",X"11",X"12",X"90",X"00",X"11",X"19",X"09",X"00",X"22",X"29",X"90",X"00",
		X"22",X"11",X"00",X"00",X"99",X"11",X"90",X"00",X"11",X"11",X"09",X"00",X"11",X"11",X"90",X"00",
		X"11",X"11",X"00",X"00",X"11",X"11",X"90",X"00",X"11",X"11",X"09",X"00",X"22",X"22",X"03",X"00",
		X"99",X"11",X"55",X"00",X"11",X"11",X"53",X"00",X"11",X"11",X"F3",X"00",X"22",X"11",X"F3",X"00",
		X"22",X"11",X"F3",X"00",X"22",X"11",X"F5",X"00",X"22",X"11",X"F3",X"00",X"22",X"22",X"F5",X"00",
		X"99",X"11",X"F5",X"00",X"11",X"11",X"F3",X"00",X"11",X"11",X"F3",X"00",X"11",X"91",X"00",X"00",
		X"19",X"E9",X"00",X"00",X"EE",X"EE",X"00",X"00",X"EE",X"EE",X"00",X"00",X"99",X"E9",X"00",X"00",
		X"22",X"FF",X"90",X"00",X"22",X"FF",X"09",X"00",X"22",X"FF",X"90",X"00",X"22",X"FF",X"00",X"00",
		X"22",X"FF",X"90",X"00",X"22",X"FF",X"09",X"00",X"29",X"FF",X"90",X"00",X"99",X"FF",X"00",X"00",
		X"22",X"FF",X"90",X"00",X"22",X"FF",X"09",X"00",X"22",X"FF",X"90",X"00",X"22",X"FF",X"00",X"00",
		X"22",X"FF",X"90",X"00",X"22",X"FF",X"09",X"00",X"32",X"FF",X"90",X"00",X"33",X"FF",X"00",X"00",
		X"33",X"FF",X"90",X"00",X"33",X"FF",X"09",X"00",X"11",X"FF",X"90",X"00",X"11",X"FF",X"00",X"00",
		X"11",X"FF",X"90",X"00",X"11",X"FF",X"09",X"00",X"11",X"FF",X"90",X"00",X"22",X"FF",X"00",X"00",
		X"11",X"FF",X"90",X"00",X"11",X"FF",X"09",X"00",X"11",X"9F",X"90",X"00",X"11",X"9F",X"00",X"00",
		X"21",X"9F",X"90",X"00",X"21",X"2F",X"09",X"00",X"21",X"9F",X"90",X"00",X"11",X"2F",X"00",X"00",
		X"99",X"39",X"00",X"00",X"EE",X"EE",X"00",X"00",X"33",X"33",X"00",X"00",X"19",X"99",X"00",X"00",
		X"11",X"91",X"00",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"22",X"22",X"F5",X"00",
		X"22",X"22",X"F5",X"00",X"99",X"92",X"F3",X"00",X"12",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",
		X"22",X"22",X"F3",X"00",X"22",X"22",X"F3",X"00",X"99",X"22",X"53",X"00",X"22",X"92",X"55",X"00",
		X"92",X"29",X"33",X"00",X"22",X"22",X"09",X"00",X"22",X"22",X"90",X"00",X"22",X"22",X"00",X"00",
		X"22",X"99",X"90",X"00",X"99",X"22",X"09",X"00",X"22",X"22",X"90",X"00",X"22",X"2F",X"00",X"00",
		X"33",X"29",X"90",X"00",X"33",X"29",X"09",X"00",X"99",X"99",X"90",X"00",X"22",X"22",X"00",X"00",
		X"22",X"29",X"90",X"00",X"22",X"29",X"09",X"00",X"22",X"29",X"90",X"00",X"22",X"29",X"00",X"00",
		X"00",X"00",X"09",X"09",X"00",X"90",X"99",X"90",X"00",X"09",X"55",X"09",X"00",X"95",X"51",X"00",
		X"09",X"55",X"51",X"99",X"00",X"55",X"11",X"99",X"09",X"55",X"11",X"55",X"95",X"55",X"11",X"33",
		X"55",X"53",X"11",X"33",X"55",X"34",X"77",X"73",X"91",X"43",X"99",X"34",X"94",X"93",X"BB",X"35",
		X"55",X"33",X"99",X"99",X"FF",X"33",X"99",X"9F",X"01",X"35",X"99",X"95",X"11",X"55",X"95",X"95",
		X"11",X"55",X"95",X"95",X"01",X"35",X"99",X"95",X"33",X"33",X"99",X"95",X"55",X"FF",X"99",X"99",
		X"94",X"FF",X"BB",X"31",X"91",X"11",X"FF",X"54",X"55",X"54",X"11",X"1F",X"F5",X"55",X"11",X"55",
		X"0F",X"55",X"11",X"55",X"00",X"55",X"11",X"FF",X"00",X"FF",X"11",X"00",X"00",X"FF",X"51",X"00",
		X"00",X"0F",X"F1",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"09",X"00",X"00",X"09",X"90",X"00",X"00",
		X"90",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"FF",X"00",X"00",
		X"F3",X"33",X"00",X"00",X"F5",X"55",X"00",X"00",X"59",X"59",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"14",X"11",X"00",X"00",X"55",X"FF",X"00",X"00",X"9F",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"09",X"00",X"00",X"09",X"90",X"00",X"00",
		X"90",X"16",X"10",X"00",X"99",X"61",X"60",X"60",X"99",X"99",X"06",X"00",X"9F",X"FF",X"00",X"00",
		X"F3",X"33",X"00",X"00",X"F5",X"55",X"00",X"00",X"59",X"59",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"14",X"11",X"00",X"00",X"55",X"FF",X"00",X"00",X"9F",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"0F",X"FF",X"66",X"00",X"00",X"00",X"10",X"00",
		X"00",X"61",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"09",X"00",X"00",X"09",X"96",X"00",X"00",
		X"90",X"69",X"00",X"00",X"99",X"99",X"00",X"00",X"99",X"99",X"60",X"00",X"9F",X"FF",X"00",X"00",
		X"F3",X"33",X"00",X"00",X"F5",X"55",X"00",X"00",X"59",X"59",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"14",X"11",X"00",X"00",X"55",X"FF",X"00",X"00",X"9F",X"09",X"00",X"00",X"90",X"90",X"00",X"00",
		X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",X"A2",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"F2",X"00",X"00",X"00",
		X"F2",X"00",X"00",X"00",X"F2",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"79",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",
		X"99",X"00",X"00",X"00",X"A9",X"90",X"00",X"00",X"DA",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"09",X"09",X"00",X"00",X"99",X"99",X"00",X"00",X"22",X"22",X"00",X"09",X"11",X"11",
		X"00",X"92",X"77",X"11",X"00",X"21",X"22",X"21",X"00",X"11",X"29",X"29",X"00",X"17",X"92",X"92",
		X"00",X"72",X"99",X"99",X"00",X"22",X"44",X"49",X"00",X"24",X"94",X"24",X"0C",X"24",X"99",X"22",
		X"C1",X"24",X"22",X"22",X"CC",X"24",X"62",X"22",X"CC",X"24",X"26",X"92",X"CC",X"24",X"92",X"22",
		X"CC",X"26",X"29",X"22",X"CC",X"24",X"92",X"22",X"CC",X"24",X"29",X"22",X"6C",X"24",X"99",X"99",
		X"CC",X"26",X"96",X"99",X"CC",X"94",X"67",X"92",X"CC",X"26",X"74",X"22",X"6C",X"94",X"44",X"24",
		X"06",X"26",X"64",X"42",X"00",X"92",X"92",X"22",X"00",X"99",X"29",X"29",X"00",X"22",X"92",X"99",
		X"00",X"11",X"99",X"92",X"00",X"17",X"22",X"21",X"00",X"01",X"11",X"11",X"00",X"00",X"71",X"20",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"92",X"09",X"00",X"00",X"11",X"99",X"09",X"00",
		X"11",X"21",X"90",X"00",X"12",X"11",X"29",X"00",X"22",X"21",X"22",X"00",X"22",X"22",X"12",X"00",
		X"99",X"22",X"11",X"00",X"77",X"22",X"21",X"00",X"72",X"99",X"22",X"00",X"27",X"26",X"92",X"00",
		X"72",X"92",X"29",X"00",X"27",X"26",X"92",X"00",X"77",X"92",X"29",X"00",X"22",X"26",X"92",X"00",
		X"22",X"92",X"29",X"00",X"22",X"26",X"92",X"00",X"22",X"92",X"29",X"00",X"22",X"26",X"92",X"00",
		X"29",X"92",X"29",X"00",X"99",X"26",X"00",X"00",X"44",X"99",X"01",X"00",X"44",X"22",X"11",X"00",
		X"44",X"92",X"11",X"00",X"22",X"29",X"10",X"00",X"92",X"99",X"00",X"00",X"99",X"12",X"00",X"00",
		X"11",X"11",X"00",X"00",X"11",X"12",X"00",X"00",X"21",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"5F",X"50",X"00",X"00",X"55",X"55",X"00",X"05",X"55",X"00",X"00",X"55",X"55",X"55",X"00",
		X"55",X"FF",X"05",X"00",X"55",X"55",X"55",X"00",X"FF",X"00",X"05",X"00",X"00",X"05",X"50",X"00",
		X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"55",X"50",X"50",X"00",X"5F",X"05",X"55",X"55",X"55",X"55",X"05",
		X"50",X"55",X"05",X"50",X"55",X"05",X"05",X"05",X"FF",X"55",X"00",X"50",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"F5",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"F5",X"00",X"00",X"00",X"5F",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"5F",X"00",X"00",X"05",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"50",X"50",X"00",X"00",X"55",X"50",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"50",X"00",X"00",X"55",X"55",X"00",X"00",
		X"5F",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"1F",X"55",X"00",X"00",
		X"15",X"15",X"50",X"00",X"11",X"11",X"55",X"00",X"11",X"11",X"55",X"00",X"F1",X"51",X"55",X"00",
		X"11",X"33",X"55",X"00",X"11",X"33",X"55",X"00",X"11",X"53",X"55",X"00",X"11",X"55",X"11",X"00",
		X"11",X"55",X"11",X"00",X"51",X"F9",X"11",X"10",X"51",X"99",X"11",X"99",X"55",X"99",X"11",X"90",
		X"55",X"9B",X"19",X"09",X"55",X"B9",X"11",X"09",X"55",X"B9",X"F1",X"99",X"55",X"B9",X"BF",X"90",
		X"55",X"BB",X"BB",X"99",X"F5",X"9B",X"9B",X"09",X"F5",X"FB",X"99",X"09",X"05",X"1F",X"9D",X"09",
		X"0F",X"91",X"DD",X"00",X"00",X"91",X"D9",X"00",X"00",X"99",X"99",X"59",X"00",X"95",X"99",X"55",
		X"99",X"99",X"12",X"99",X"99",X"99",X"91",X"99",X"99",X"19",X"99",X"99",X"99",X"12",X"93",X"F9",
		X"99",X"55",X"FF",X"00",X"90",X"55",X"99",X"99",X"90",X"00",X"9F",X"99",X"00",X"99",X"F9",X"FF",
		X"90",X"99",X"99",X"00",X"09",X"00",X"9F",X"F0",X"00",X"09",X"F9",X"F0",X"00",X"09",X"39",X"1F",
		X"00",X"00",X"19",X"11",X"00",X"00",X"12",X"99",X"00",X"00",X"F1",X"90",X"00",X"00",X"F1",X"99",
		X"00",X"00",X"9F",X"09",X"00",X"00",X"9F",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"99",X"09",X"DD",X"00",X"00",X"05",X"BB",X"00",X"00",X"09",X"99",
		X"00",X"99",X"00",X"99",X"00",X"BA",X"99",X"99",X"00",X"AB",X"D9",X"99",X"09",X"4A",X"9D",X"99",
		X"9D",X"B4",X"D9",X"99",X"DD",X"99",X"99",X"99",X"DD",X"94",X"BA",X"BB",X"DD",X"4F",X"BB",X"BB",
		X"99",X"FF",X"BB",X"B9",X"9B",X"FF",X"BB",X"B5",X"9B",X"FF",X"BB",X"B9",X"9B",X"FF",X"BB",X"BF",
		X"9B",X"F9",X"BB",X"59",X"9F",X"FF",X"FB",X"B5",X"9A",X"99",X"BF",X"B9",X"BB",X"49",X"FB",X"B5",
		X"BB",X"F4",X"FB",X"BB",X"BB",X"F9",X"99",X"99",X"AB",X"94",X"AA",X"99",X"0A",X"4B",X"AA",X"99",
		X"00",X"BB",X"99",X"99",X"00",X"BB",X"90",X"99",X"00",X"99",X"00",X"99",X"00",X"00",X"09",X"99",
		X"00",X"00",X"05",X"DD",X"00",X"99",X"09",X"BB",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",
		X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",
		X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"A0",X"D9",X"A9",X"00",X"A0",
		X"DB",X"DB",X"E0",X"A0",X"BD",X"BD",X"D9",X"90",X"BB",X"BB",X"BB",X"AA",X"FF",X"FF",X"FF",X"FF",
		X"55",X"55",X"BB",X"AA",X"BB",X"BB",X"BA",X"A0",X"DB",X"DB",X"E0",X"B0",X"DD",X"AA",X"00",X"A0",
		X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",X"A0",
		X"00",X"00",X"00",X"BA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"99",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",X"00",X"D4",X"00",X"00",
		X"02",X"94",X"90",X"00",X"02",X"BB",X"D9",X"00",X"02",X"B4",X"DD",X"90",X"99",X"B4",X"DD",X"99",
		X"AB",X"4F",X"AD",X"D9",X"0A",X"4F",X"BA",X"DD",X"0A",X"9F",X"BA",X"DD",X"09",X"FF",X"BB",X"9B",
		X"09",X"99",X"BB",X"99",X"00",X"9F",X"BB",X"99",X"00",X"49",X"BB",X"99",X"00",X"49",X"BB",X"99",
		X"00",X"F4",X"BB",X"99",X"00",X"44",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"90",X"BB",X"BB",X"99",
		X"99",X"AA",X"BB",X"B9",X"00",X"9A",X"BF",X"FB",X"00",X"09",X"99",X"9B",X"00",X"09",X"99",X"BB",
		X"00",X"99",X"90",X"FB",X"00",X"90",X"E0",X"B9",X"00",X"99",X"09",X"99",X"00",X"09",X"99",X"9D",
		X"00",X"00",X"99",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"B9",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"BD",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"BF",X"D0",X"00",X"00",X"BB",X"DD",X"00",X"00",X"DB",X"BB",X"00",X"00",
		X"DD",X"BB",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",
		X"00",X"BB",X"00",X"D0",X"00",X"DD",X"D0",X"D0",X"00",X"00",X"BD",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"BD",X"00",
		X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",
		X"00",X"00",X"B0",X"00",X"00",X"00",X"BB",X"B0",X"00",X"00",X"AA",X"B0",X"00",X"00",X"A0",X"B0",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"49",X"00",X"00",X"2F",X"49",X"00",X"00",X"FB",X"44",X"00",X"00",X"BB",X"F4",X"90",X"00",
		X"FB",X"94",X"90",X"00",X"BB",X"F4",X"99",X"00",X"F4",X"94",X"99",X"00",X"44",X"94",X"09",X"00",
		X"F4",X"44",X"00",X"00",X"F4",X"44",X"00",X"00",X"F4",X"4B",X"99",X"00",X"F4",X"BB",X"90",X"00",
		X"94",X"BB",X"90",X"00",X"94",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",X"44",X"BB",X"00",X"00",
		X"B9",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"AA",X"BB",X"00",X"00",X"AA",X"BB",X"09",X"00",
		X"AA",X"BB",X"99",X"00",X"AA",X"BB",X"99",X"90",X"09",X"BB",X"99",X"90",X"00",X"B9",X"99",X"00",
		X"09",X"99",X"99",X"00",X"09",X"9B",X"90",X"00",X"90",X"0B",X"E0",X"00",X"90",X"9B",X"A0",X"00",
		X"00",X"9B",X"A0",X"00",X"90",X"99",X"A0",X"00",X"00",X"99",X"BA",X"00",X"D0",X"90",X"BD",X"00",
		X"DD",X"00",X"BD",X"00",X"BD",X"00",X"5B",X"00",X"BB",X"00",X"FB",X"00",X"0B",X"00",X"FB",X"00",
		X"00",X"00",X"B5",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"DB",X"00",
		X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",
		X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",X"00",X"00",X"D0",X"00",X"00",X"A0",X"DA",
		X"00",X"00",X"A0",X"BD",X"00",X"00",X"AA",X"BA",X"00",X"00",X"9A",X"DA",X"00",X"00",X"09",X"0D",
		X"BD",X"BB",X"B0",X"D9",X"BD",X"09",X"00",X"D9",X"0D",X"09",X"00",X"D0",X"00",X"0D",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",
		X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"0D",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"BF",X"AA",X"00",X"00",X"BB",X"AA",X"00",X"00",X"BB",X"AA",X"00",
		X"00",X"AB",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"A2",X"A0",X"00",X"00",X"AA",X"A0",X"00",X"00",X"BB",X"D9",X"00",X"00",X"BB",X"DD",X"00",
		X"00",X"BB",X"DD",X"00",X"00",X"BA",X"DD",X"00",X"09",X"AA",X"9D",X"00",X"09",X"AA",X"99",X"00",
		X"09",X"4B",X"44",X"00",X"09",X"F4",X"9B",X"00",X"09",X"FF",X"9B",X"00",X"09",X"F4",X"9B",X"00",
		X"09",X"F4",X"99",X"00",X"09",X"94",X"94",X"00",X"09",X"49",X"49",X"00",X"09",X"44",X"49",X"00",
		X"09",X"FB",X"F9",X"00",X"09",X"BF",X"B9",X"00",X"00",X"9B",X"99",X"00",X"00",X"9F",X"9D",X"00",
		X"00",X"9B",X"9D",X"00",X"90",X"9F",X"9D",X"95",X"90",X"9A",X"9D",X"99",X"9D",X"9F",X"9D",X"D9",
		X"BD",X"9A",X"99",X"D9",X"BD",X"9B",X"99",X"D9",X"BD",X"99",X"90",X"D9",X"BD",X"99",X"99",X"D9",
		X"BD",X"BB",X"B9",X"D9",X"BD",X"59",X"B9",X"D9",X"BD",X"B9",X"B9",X"D9",X"BD",X"59",X"B9",X"D9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D0",
		X"00",X"00",X"00",X"D0",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"DD",X"00",X"00",X"00",X"0D",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",
		X"00",X"00",X"99",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"46",X"00",
		X"00",X"00",X"60",X"00",X"00",X"00",X"40",X"00",X"00",X"40",X"00",X"00",X"00",X"64",X"44",X"00",
		X"00",X"66",X"66",X"00",X"00",X"06",X"66",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"40",X"06",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"40",X"00",X"00",X"60",X"66",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"46",X"00",X"00",X"04",X"66",X"00",X"00",X"46",X"46",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"66",X"00",X"00",X"00",X"66",X"40",
		X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"46",X"00",X"00",X"00",X"66",X"00",
		X"44",X"00",X"60",X"00",X"06",X"00",X"40",X"00",X"00",X"40",X"60",X"00",X"00",X"64",X"66",X"00",
		X"00",X"66",X"64",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"40",X"60",X"66",X"00",X"66",X"00",X"06",X"00",X"66",X"00",X"04",X"00",
		X"00",X"00",X"40",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"06",X"00",
		X"00",X"00",X"66",X"00",X"00",X"66",X"46",X"00",X"00",X"64",X"66",X"00",X"00",X"46",X"46",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"66",X"00",X"06",X"00",X"66",X"00",
		X"00",X"00",X"66",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",
		X"00",X"04",X"00",X"00",X"06",X"66",X"00",X"00",X"00",X"60",X"46",X"00",X"00",X"06",X"66",X"00",
		X"44",X"04",X"60",X"00",X"46",X"00",X"40",X"00",X"66",X"40",X"60",X"00",X"60",X"00",X"66",X"00",
		X"00",X"04",X"64",X"00",X"00",X"46",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"64",X"00",
		X"64",X"00",X"66",X"00",X"66",X"60",X"66",X"00",X"66",X"44",X"06",X"00",X"66",X"66",X"04",X"00",
		X"00",X"66",X"40",X"00",X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"66",X"00",
		X"00",X"06",X"44",X"60",X"64",X"66",X"66",X"00",X"66",X"64",X"66",X"00",X"06",X"66",X"46",X"00",
		X"00",X"66",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"60",X"66",X"00",X"66",X"00",X"66",X"00",
		X"04",X"40",X"66",X"00",X"00",X"66",X"04",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"46",X"06",X"00",X"00",X"66",X"60",
		X"44",X"00",X"60",X"60",X"46",X"00",X"40",X"00",X"66",X"40",X"60",X"00",X"66",X"00",X"66",X"00",
		X"06",X"04",X"64",X"00",X"00",X"46",X"66",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"64",X"40",
		X"60",X"00",X"66",X"66",X"60",X"00",X"66",X"00",X"00",X"40",X"06",X"00",X"00",X"00",X"04",X"00",
		X"00",X"00",X"40",X"00",X"06",X"60",X"66",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"66",X"06",
		X"00",X"00",X"44",X"60",X"64",X"40",X"66",X"00",X"40",X"00",X"66",X"00",X"46",X"06",X"46",X"00",
		X"66",X"00",X"66",X"00",X"60",X"00",X"66",X"00",X"00",X"00",X"66",X"60",X"00",X"00",X"66",X"06",
		X"04",X"40",X"66",X"00",X"00",X"6E",X"04",X"00",X"00",X"EE",X"00",X"40",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",
		X"00",X"00",X"00",X"00",X"00",X"A0",X"A0",X"00",X"00",X"00",X"0A",X"0A",X"00",X"0A",X"A0",X"00",
		X"0A",X"A0",X"0A",X"00",X"00",X"0A",X"AF",X"00",X"A0",X"00",X"F0",X"00",X"0A",X"0A",X"00",X"00",
		X"00",X"F0",X"0F",X"00",X"AF",X"0F",X"00",X"F0",X"0F",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"0A",X"A0",X"00",X"00",X"A0",X"00",X"00",X"00",
		X"F0",X"0A",X"0A",X"00",X"0F",X"A0",X"A0",X"00",X"F0",X"00",X"0A",X"0A",X"0F",X"FF",X"A0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"0A",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"0A",X"00",X"00",X"A0",X"00",
		X"0A",X"0A",X"0F",X"00",X"A0",X"0F",X"F0",X"00",X"0A",X"F0",X"0F",X"F0",X"F0",X"0F",X"00",X"00",
		X"0A",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"FA",X"A0",X"00",X"00",X"00",X"00",X"A0",X"00",
		X"0F",X"FA",X"0A",X"00",X"F0",X"0F",X"A0",X"00",X"00",X"00",X"0F",X"0A",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"F0",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"FF",X"F0",X"00",X"FF",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"0F",X"FF",X"00",X"00",X"00",X"F0",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"0F",X"F0",X"00",
		X"FF",X"F0",X"0F",X"00",X"FF",X"0F",X"FF",X"00",X"00",X"F0",X"F0",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"F0",X"FF",X"00",X"00",X"FF",X"0F",X"00",X"F0",X"F0",X"FF",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"FF",X"FF",X"00",X"00",X"FF",X"FF",X"F0",X"00",X"F0",X"0F",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"0F",X"F0",X"FF",X"F0",X"0F",X"00",X"F0",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"0F",X"0F",X"00",
		X"00",X"F0",X"F0",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"FF",X"F0",X"F0",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",
		X"0F",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"B3",X"93",X"00",X"09",X"5B",X"BB",X"00",
		X"09",X"5F",X"BB",X"00",X"00",X"B3",X"93",X"00",X"00",X"39",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"39",X"00",X"00",X"00",X"B3",X"93",X"00",X"09",X"55",X"BB",X"00",
		X"09",X"5F",X"BB",X"00",X"00",X"B3",X"93",X"00",X"00",X"39",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"93",X"00",X"00",X"30",X"30",X"09",X"00",X"50",X"00",X"00",X"05",
		X"05",X"05",X"05",X"00",X"30",X"30",X"5F",X"50",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"00",X"0F",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"93",X"93",X"00",X"00",X"30",X"30",X"09",X"00",X"50",X"00",X"00",X"00",
		X"05",X"05",X"05",X"0F",X"30",X"30",X"50",X"50",X"03",X"03",X"03",X"00",X"00",X"00",X"00",X"00",
		X"05",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"05",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"09",X"99",X"99",X"00",X"9D",X"99",X"99",
		X"00",X"DD",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"DD",X"99",X"99",X"00",X"99",X"99",X"99",
		X"09",X"DE",X"EE",X"55",X"9D",X"99",X"B5",X"99",X"DD",X"DE",X"5B",X"EE",X"99",X"EE",X"B5",X"99",
		X"DD",X"E9",X"99",X"AB",X"99",X"E9",X"FE",X"BA",X"DD",X"99",X"F9",X"AB",X"99",X"EE",X"F5",X"BA",
		X"AA",X"BB",X"F5",X"AB",X"AB",X"99",X"F9",X"BA",X"BA",X"59",X"F5",X"AB",X"AB",X"B9",X"B5",X"9A",
		X"BA",X"5B",X"5B",X"99",X"AB",X"A5",X"55",X"FF",X"BA",X"BB",X"5B",X"99",X"0B",X"A5",X"55",X"55",
		X"00",X"BA",X"99",X"95",X"00",X"AB",X"99",X"99",X"00",X"BA",X"BA",X"AA",X"00",X"AB",X"AB",X"BB",
		X"00",X"BA",X"BA",X"AA",X"00",X"BB",X"AB",X"BB",X"00",X"00",X"BA",X"BA",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"99",X"9D",X"9D",X"00",
		X"99",X"DD",X"99",X"00",X"99",X"9D",X"99",X"00",X"9E",X"BB",X"99",X"00",X"99",X"DD",X"99",X"00",
		X"EE",X"BB",X"99",X"00",X"9E",X"DD",X"99",X"00",X"E9",X"BB",X"99",X"00",X"AE",X"DD",X"99",X"00",
		X"E9",X"BB",X"99",X"00",X"A9",X"BB",X"99",X"00",X"99",X"BB",X"99",X"00",X"A9",X"BB",X"99",X"00",
		X"99",X"AB",X"99",X"00",X"A9",X"BB",X"99",X"00",X"99",X"AB",X"99",X"00",X"A9",X"BB",X"99",X"00",
		X"99",X"AA",X"99",X"00",X"99",X"BB",X"99",X"00",X"99",X"AA",X"99",X"00",X"99",X"BB",X"99",X"00",
		X"59",X"AA",X"99",X"00",X"55",X"BB",X"99",X"00",X"AA",X"AA",X"A9",X"00",X"BA",X"BA",X"AA",X"00",
		X"AA",X"AA",X"AA",X"00",X"AB",X"AA",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"9A",X"9A",X"00",X"AB",X"AB",X"AB",X"00",X"BD",X"BD",X"BD",X"00",X"BB",X"BB",X"BB",
		X"00",X"5B",X"5B",X"5B",X"00",X"BA",X"BA",X"BA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"99",X"00",X"BA",X"BA",X"BA",
		X"00",X"AB",X"AB",X"AB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"AB",X"AB",X"AB",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"0F",X"00",X"0F",X"F0",X"0F",X"00",X"FF",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"F0",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"0F",X"00",X"00",X"F5",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"F0",X"00",X"00",X"0F",X"0F",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"F0",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"0F",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"0F",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"05",X"0F",X"00",X"00",X"00",X"00",X"0F",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"0F",X"00",
		X"00",X"0F",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"F0",X"FF",X"0F",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",
		X"0F",X"FF",X"00",X"00",X"F0",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"F0",X"00",
		X"00",X"0F",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"F0",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"5F",X"0F",X"00",X"00",X"50",X"00",X"00",X"F0",X"0F",X"00",
		X"00",X"0F",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",
		X"00",X"00",X"05",X"05",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"FA",X"00",X"00",X"00",X"A5",X"A0",X"00",X"99",X"99",X"00",X"00",X"95",X"55",X"0F",
		X"00",X"99",X"55",X"99",X"00",X"99",X"55",X"55",X"00",X"95",X"55",X"33",X"09",X"55",X"11",X"33",
		X"00",X"33",X"77",X"77",X"00",X"44",X"33",X"99",X"00",X"77",X"3A",X"B3",X"08",X"13",X"AB",X"99",
		X"00",X"55",X"BB",X"99",X"88",X"55",X"B9",X"9D",X"00",X"53",X"B9",X"9D",X"00",X"F5",X"B9",X"9D",
		X"00",X"FF",X"B9",X"9D",X"80",X"FF",X"BB",X"99",X"00",X"9F",X"A9",X"99",X"00",X"19",X"99",X"B3",
		X"08",X"11",X"F9",X"FF",X"99",X"55",X"11",X"11",X"00",X"99",X"11",X"55",X"00",X"59",X"55",X"55",
		X"00",X"99",X"55",X"5F",X"00",X"08",X"55",X"90",X"00",X"09",X"F5",X"90",X"00",X"00",X"99",X"90",
		X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"90",X"09",X"30",X"00",X"59",X"99",X"03",X"00",
		X"5F",X"9F",X"30",X"00",X"95",X"33",X"03",X"00",X"11",X"11",X"30",X"00",X"99",X"99",X"00",X"00",
		X"9F",X"FF",X"00",X"00",X"9F",X"60",X"00",X"00",X"9F",X"F0",X"00",X"00",X"9F",X"FF",X"00",X"00",
		X"9F",X"9F",X"00",X"00",X"9F",X"FF",X"F0",X"00",X"99",X"99",X"F0",X"00",X"41",X"11",X"F0",X"00",
		X"55",X"FF",X"00",X"00",X"F9",X"99",X"00",X"00",X"FF",X"99",X"00",X"00",X"00",X"F9",X"00",X"00",
		X"0F",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"F0",X"00",X"00",
		X"0F",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"0F",X"00",X"0F",X"0F",X"0F",X"00",X"09",X"00",X"00",X"00",X"90",X"55",X"00",
		X"00",X"59",X"59",X"00",X"00",X"95",X"55",X"35",X"00",X"55",X"55",X"53",X"00",X"55",X"31",X"33",
		X"00",X"93",X"77",X"77",X"00",X"14",X"33",X"99",X"00",X"47",X"33",X"BB",X"00",X"71",X"3A",X"99",
		X"00",X"55",X"AB",X"99",X"08",X"55",X"AB",X"99",X"00",X"55",X"AB",X"99",X"00",X"FF",X"AB",X"99",
		X"00",X"FF",X"AB",X"99",X"08",X"FF",X"AB",X"99",X"00",X"11",X"99",X"99",X"00",X"41",X"99",X"99",
		X"00",X"11",X"99",X"99",X"99",X"55",X"19",X"99",X"00",X"55",X"59",X"95",X"00",X"99",X"59",X"55",
		X"00",X"99",X"59",X"00",X"00",X"00",X"59",X"00",X"00",X"00",X"F9",X"00",X"00",X"00",X"99",X"99",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"FF",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"F0",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"50",X"00",X"03",X"00",X"55",X"00",X"30",X"00",
		X"95",X"00",X"03",X"00",X"99",X"00",X"30",X"00",X"11",X"F0",X"03",X"00",X"99",X"F0",X"00",X"00",
		X"99",X"F0",X"F0",X"00",X"59",X"00",X"00",X"0F",X"59",X"0F",X"00",X"00",X"59",X"00",X"00",X"0F",
		X"59",X"00",X"F0",X"0F",X"99",X"00",X"0F",X"0F",X"99",X"90",X"00",X"00",X"44",X"10",X"0F",X"00",
		X"55",X"F0",X"F0",X"00",X"FF",X"90",X"F0",X"00",X"FF",X"F0",X"00",X"00",X"00",X"0F",X"F0",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",X"F0",X"00",X"0F",X"0F",X"00",X"00",
		X"00",X"00",X"0F",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"F0",X"00",X"F0",X"F0",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",X"0F",X"0F",X"0F",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"55",X"00",X"F0",X"55",X"55",X"53",
		X"00",X"55",X"31",X"33",X"0F",X"53",X"77",X"77",X"F0",X"14",X"33",X"99",X"00",X"47",X"33",X"00",
		X"00",X"71",X"3A",X"00",X"00",X"55",X"AB",X"00",X"08",X"55",X"AB",X"00",X"00",X"55",X"9B",X"00",
		X"00",X"FF",X"9B",X"00",X"00",X"FF",X"9B",X"99",X"08",X"FF",X"9B",X"99",X"00",X"99",X"9A",X"99",
		X"00",X"49",X"99",X"99",X"00",X"11",X"99",X"99",X"99",X"55",X"19",X"99",X"00",X"95",X"55",X"11",
		X"00",X"99",X"55",X"15",X"00",X"99",X"55",X"15",X"00",X"00",X"55",X"55",X"00",X"00",X"99",X"99",
		X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"03",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"F0",X"00",X"F0",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"99",X"00",X"0F",X"00",X"99",X"00",X"00",X"00",
		X"44",X"00",X"0F",X"00",X"55",X"0F",X"F0",X"00",X"FF",X"0F",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"0F",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"F0",X"00",X"FF",X"F0",X"0F",X"00",X"FF",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"0F",X"09",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",
		X"00",X"00",X"33",X"00",X"00",X"05",X"47",X"00",X"00",X"99",X"93",X"00",X"00",X"44",X"33",X"0B",
		X"00",X"55",X"33",X"00",X"00",X"11",X"55",X"00",X"00",X"95",X"55",X"00",X"0F",X"55",X"5A",X"00",
		X"00",X"9F",X"90",X"00",X"00",X"9F",X"99",X"09",X"00",X"11",X"99",X"00",X"00",X"55",X"99",X"09",
		X"0F",X"44",X"9F",X"90",X"00",X"10",X"99",X"FF",X"00",X"05",X"41",X"19",X"00",X"00",X"55",X"F9",
		X"00",X"09",X"55",X"F0",X"00",X"00",X"55",X"09",X"00",X"F0",X"00",X"99",X"F0",X"0F",X"00",X"00",
		X"0F",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"00",X"F0",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"F0",X"0F",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"F0",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"F0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"51",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"0F",X"00",X"F0",X"00",X"F0",X"00",X"00",X"0F",X"00",X"00",X"0F",X"F0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",
		X"00",X"39",X"90",X"00",X"99",X"33",X"90",X"00",X"91",X"FF",X"90",X"00",X"91",X"55",X"99",X"90",
		X"51",X"F5",X"F9",X"00",X"55",X"55",X"F9",X"90",X"55",X"11",X"59",X"90",X"55",X"11",X"55",X"90",
		X"F5",X"99",X"51",X"99",X"F5",X"99",X"11",X"90",X"FF",X"5F",X"11",X"90",X"FF",X"55",X"11",X"09",
		X"1F",X"FF",X"91",X"90",X"99",X"F9",X"99",X"39",X"99",X"F9",X"BF",X"33",X"99",X"F9",X"9B",X"F3",
		X"99",X"F9",X"99",X"F3",X"59",X"F9",X"99",X"59",X"50",X"FB",X"99",X"5F",X"90",X"1F",X"99",X"5F",
		X"99",X"11",X"99",X"99",X"99",X"11",X"99",X"F9",X"99",X"11",X"99",X"99",X"99",X"51",X"1F",X"99",
		X"09",X"52",X"11",X"99",X"00",X"55",X"51",X"00",X"00",X"55",X"55",X"99",X"00",X"F5",X"5F",X"99",
		X"00",X"F5",X"FF",X"9F",X"00",X"FF",X"0F",X"FF",X"00",X"FF",X"00",X"FF",X"00",X"0F",X"00",X"FF",
		X"F0",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"9F",X"11",X"00",X"00",X"99",X"11",X"99",X"00",
		X"99",X"11",X"FF",X"00",X"00",X"00",X"F0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"90",X"00",X"00",X"00",X"99",X"00",X"09",X"00",X"09",X"00",X"99",X"00",X"09",X"99",X"9F",X"00",
		X"09",X"FF",X"F5",X"00",X"00",X"59",X"55",X"00",X"00",X"11",X"11",X"00",X"00",X"11",X"99",X"00",
		X"00",X"FF",X"FF",X"00",X"09",X"F9",X"FF",X"00",X"90",X"F9",X"FF",X"00",X"09",X"F9",X"FF",X"00",
		X"99",X"F9",X"FF",X"00",X"9F",X"FF",X"FF",X"00",X"F9",X"99",X"99",X"00",X"00",X"11",X"11",X"00",
		X"00",X"11",X"1F",X"00",X"09",X"99",X"9F",X"00",X"99",X"99",X"99",X"00",X"09",X"0F",X"99",X"00",
		X"00",X"00",X"F9",X"00",X"00",X"00",X"0F",X"00",X"00",X"90",X"00",X"00",X"09",X"99",X"00",X"00",
		X"92",X"99",X"99",X"99",X"29",X"22",X"22",X"22",X"92",X"22",X"22",X"92",X"99",X"99",X"99",X"99",
		X"CC",X"22",X"22",X"22",X"C9",X"22",X"22",X"22",X"9C",X"92",X"22",X"22",X"9C",X"C9",X"99",X"99",
		X"99",X"29",X"C2",X"22",X"29",X"99",X"22",X"22",X"22",X"99",X"92",X"22",X"22",X"22",X"9C",X"99",
		X"22",X"22",X"C9",X"99",X"22",X"22",X"22",X"29",X"99",X"C2",X"22",X"22",X"93",X"99",X"22",X"29",
		X"93",X"99",X"9C",X"99",X"93",X"22",X"C9",X"C2",X"93",X"22",X"22",X"22",X"93",X"22",X"22",X"2C",
		X"99",X"C9",X"92",X"22",X"00",X"C2",X"99",X"99",X"02",X"CC",X"22",X"29",X"02",X"2C",X"22",X"22",
		X"03",X"22",X"22",X"CC",X"99",X"92",X"9C",X"99",X"CC",X"99",X"29",X"99",X"92",X"22",X"22",X"C3",
		X"CC",X"22",X"C2",X"33",X"3C",X"C2",X"22",X"33",X"3C",X"2C",X"22",X"99",X"9C",X"22",X"22",X"33",
		X"99",X"99",X"99",X"F0",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"00",X"99",X"99",X"99",X"F0",
		X"22",X"22",X"22",X"2F",X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"00",X"99",X"99",X"99",X"90",
		X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"F2",X"22",X"92",X"99",X"00",X"99",X"99",X"99",X"FF",
		X"00",X"00",X"F0",X"20",X"99",X"00",X"FF",X"00",X"92",X"99",X"00",X"FF",X"99",X"92",X"F0",X"F0",
		X"22",X"22",X"FF",X"0F",X"99",X"99",X"F0",X"F0",X"92",X"92",X"F0",X"00",X"22",X"29",X"00",X"00",
		X"22",X"92",X"2F",X"F0",X"99",X"22",X"0F",X"00",X"99",X"99",X"FF",X"00",X"C9",X"92",X"00",X"00",
		X"C2",X"22",X"F0",X"0F",X"22",X"92",X"0F",X"F0",X"39",X"22",X"00",X"F0",X"99",X"99",X"F0",X"0F",
		X"92",X"29",X"0F",X"F0",X"92",X"22",X"00",X"00",X"92",X"92",X"20",X"00",X"92",X"22",X"0F",X"00",
		X"29",X"99",X"99",X"99",X"20",X"22",X"22",X"22",X"22",X"C2",X"22",X"22",X"22",X"C2",X"22",X"2C",
		X"C2",X"99",X"92",X"99",X"C9",X"99",X"92",X"22",X"C2",X"22",X"09",X"22",X"CC",X"22",X"90",X"22",
		X"3C",X"22",X"09",X"22",X"9C",X"22",X"90",X"22",X"C9",X"99",X"99",X"92",X"C2",X"22",X"29",X"22",
		X"CC",X"22",X"22",X"92",X"0C",X"22",X"22",X"22",X"02",X"22",X"22",X"22",X"02",X"99",X"99",X"9C",
		X"9C",X"99",X"29",X"29",X"33",X"22",X"22",X"22",X"33",X"22",X"C2",X"22",X"33",X"2C",X"C2",X"92",
		X"99",X"C2",X"22",X"99",X"33",X"CC",X"99",X"00",X"99",X"90",X"0F",X"00",X"99",X"29",X"F0",X"00",
		X"99",X"22",X"F0",X"00",X"99",X"22",X"00",X"00",X"09",X"99",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F0",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"00",X"0F",X"00",X"00",X"0F",X"FF",X"00",X"00",
		X"39",X"99",X"00",X"F0",X"29",X"22",X"00",X"00",X"22",X"92",X"2F",X"00",X"29",X"22",X"00",X"00",
		X"22",X"29",X"0F",X"F0",X"39",X"32",X"0F",X"00",X"92",X"92",X"00",X"00",X"22",X"22",X"00",X"FF",
		X"29",X"92",X"20",X"0F",X"99",X"22",X"0F",X"00",X"22",X"99",X"00",X"0F",X"22",X"22",X"0F",X"00",
		X"22",X"29",X"00",X"0F",X"92",X"22",X"00",X"00",X"99",X"92",X"02",X"00",X"22",X"22",X"0F",X"00",
		X"22",X"29",X"0F",X"00",X"29",X"92",X"0F",X"00",X"22",X"99",X"00",X"00",X"99",X"00",X"F0",X"00",
		X"0F",X"00",X"00",X"0F",X"00",X"FF",X"F0",X"0F",X"0F",X"F0",X"2F",X"00",X"0F",X"F2",X"00",X"00",
		X"00",X"29",X"0F",X"00",X"00",X"92",X"20",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"00",X"0F",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"0F",X"00",
		X"92",X"99",X"99",X"99",X"29",X"22",X"22",X"22",X"92",X"22",X"22",X"92",X"99",X"99",X"99",X"99",
		X"CC",X"22",X"22",X"22",X"C9",X"22",X"22",X"22",X"9C",X"92",X"22",X"22",X"9C",X"C9",X"99",X"99",
		X"99",X"29",X"C2",X"22",X"29",X"99",X"22",X"22",X"22",X"99",X"92",X"22",X"22",X"22",X"9C",X"99",
		X"22",X"22",X"C9",X"99",X"22",X"22",X"22",X"29",X"99",X"C2",X"22",X"22",X"93",X"99",X"22",X"29",
		X"93",X"99",X"9C",X"99",X"93",X"22",X"C9",X"C2",X"93",X"22",X"22",X"22",X"93",X"22",X"22",X"2C",
		X"99",X"C9",X"92",X"22",X"00",X"C2",X"99",X"99",X"02",X"CC",X"22",X"29",X"02",X"2C",X"22",X"22",
		X"03",X"22",X"22",X"CC",X"99",X"92",X"9C",X"99",X"CC",X"99",X"29",X"99",X"92",X"22",X"22",X"C3",
		X"CC",X"22",X"C2",X"33",X"3C",X"C2",X"22",X"33",X"3C",X"2C",X"22",X"99",X"9C",X"22",X"22",X"33",
		X"99",X"99",X"99",X"00",X"22",X"22",X"22",X"00",X"22",X"22",X"22",X"F0",X"99",X"99",X"99",X"0F",
		X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"00",X"99",X"99",X"99",X"90",
		X"22",X"22",X"22",X"20",X"22",X"22",X"22",X"92",X"22",X"92",X"99",X"00",X"99",X"99",X"99",X"00",
		X"00",X"00",X"00",X"20",X"99",X"00",X"00",X"00",X"92",X"99",X"00",X"FF",X"99",X"92",X"00",X"00",
		X"22",X"22",X"00",X"00",X"99",X"99",X"20",X"00",X"92",X"92",X"00",X"00",X"22",X"29",X"00",X"00",
		X"22",X"92",X"20",X"F0",X"99",X"22",X"00",X"0F",X"99",X"99",X"00",X"F0",X"C9",X"92",X"00",X"0F",
		X"C2",X"22",X"0F",X"0F",X"22",X"92",X"00",X"F0",X"39",X"22",X"F0",X"00",X"99",X"99",X"20",X"00",
		X"92",X"29",X"F0",X"F0",X"92",X"22",X"F0",X"00",X"92",X"92",X"20",X"F0",X"92",X"22",X"00",X"00",
		X"29",X"99",X"99",X"99",X"20",X"22",X"22",X"22",X"22",X"C2",X"22",X"22",X"22",X"C2",X"22",X"2C",
		X"C2",X"99",X"92",X"99",X"C9",X"99",X"92",X"22",X"C2",X"22",X"09",X"22",X"CC",X"22",X"90",X"22",
		X"3C",X"22",X"09",X"22",X"9C",X"22",X"90",X"22",X"C9",X"99",X"99",X"92",X"C2",X"22",X"29",X"22",
		X"CC",X"22",X"22",X"92",X"0C",X"22",X"22",X"22",X"02",X"22",X"22",X"22",X"02",X"99",X"99",X"9C",
		X"9C",X"99",X"29",X"29",X"33",X"22",X"22",X"22",X"33",X"22",X"C2",X"22",X"33",X"2C",X"C2",X"92",
		X"99",X"C2",X"22",X"99",X"33",X"CC",X"99",X"00",X"99",X"90",X"F0",X"00",X"99",X"29",X"F0",X"00",
		X"99",X"22",X"00",X"00",X"99",X"22",X"00",X"00",X"09",X"99",X"F0",X"00",X"00",X"00",X"0F",X"00",
		X"00",X"00",X"F0",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",
		X"39",X"99",X"9F",X"00",X"29",X"22",X"00",X"0F",X"22",X"92",X"2F",X"00",X"29",X"22",X"00",X"F0",
		X"22",X"29",X"0F",X"F0",X"39",X"32",X"02",X"F0",X"92",X"92",X"00",X"F0",X"22",X"22",X"00",X"00",
		X"29",X"92",X"20",X"FF",X"99",X"22",X"00",X"0F",X"22",X"99",X"00",X"00",X"22",X"22",X"00",X"0F",
		X"22",X"29",X"00",X"F0",X"92",X"22",X"0F",X"0F",X"99",X"92",X"02",X"0F",X"22",X"22",X"0F",X"0F",
		X"22",X"29",X"00",X"F0",X"29",X"92",X"0F",X"00",X"22",X"99",X"00",X"00",X"99",X"0F",X"F0",X"00",
		X"00",X"F0",X"00",X"00",X"00",X"00",X"F0",X"F0",X"00",X"F0",X"20",X"F0",X"00",X"F2",X"00",X"00",
		X"00",X"29",X"00",X"00",X"00",X"92",X"20",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",
		X"00",X"99",X"0F",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",X"00",X"99",X"F0",X"00",
		X"0F",X"A0",X"00",X"00",X"0F",X"AA",X"00",X"00",X"FF",X"E9",X"00",X"00",X"FF",X"E7",X"AA",X"00",
		X"F0",X"EA",X"99",X"00",X"F0",X"EE",X"99",X"AA",X"FF",X"EE",X"99",X"99",X"F3",X"55",X"99",X"99",
		X"09",X"99",X"3A",X"99",X"59",X"93",X"53",X"A3",X"59",X"3A",X"7A",X"33",X"59",X"AA",X"AA",X"F9",
		X"59",X"AF",X"AA",X"59",X"59",X"FF",X"99",X"59",X"59",X"FF",X"99",X"59",X"59",X"FF",X"55",X"59",
		X"9F",X"FF",X"A5",X"99",X"99",X"EF",X"AA",X"99",X"A3",X"EE",X"AA",X"99",X"9A",X"EE",X"AA",X"99",
		X"93",X"99",X"AA",X"9E",X"93",X"E9",X"EE",X"99",X"99",X"AE",X"E5",X"99",X"59",X"EE",X"9E",X"99",
		X"D9",X"AE",X"9E",X"99",X"09",X"EA",X"99",X"99",X"0D",X"5A",X"99",X"99",X"00",X"D9",X"99",X"FF",
		X"00",X"00",X"99",X"99",X"00",X"00",X"D9",X"99",X"00",X"00",X"00",X"D9",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"09",X"00",X"00",X"99",X"99",X"90",X"00",
		X"99",X"3A",X"00",X"00",X"99",X"99",X"99",X"00",X"A9",X"99",X"99",X"00",X"AA",X"99",X"99",X"00",
		X"AA",X"A7",X"99",X"F0",X"AA",X"AA",X"9A",X"F0",X"AA",X"AA",X"99",X"F0",X"AA",X"94",X"99",X"F0",
		X"AA",X"AA",X"99",X"00",X"AA",X"AA",X"F9",X"00",X"AA",X"AA",X"F9",X"00",X"AA",X"9A",X"F9",X"00",
		X"AA",X"AA",X"F9",X"00",X"AA",X"9A",X"F9",X"00",X"AA",X"AA",X"F9",X"00",X"AE",X"AA",X"F9",X"00",
		X"AE",X"AA",X"99",X"00",X"EE",X"AA",X"99",X"00",X"EE",X"AA",X"99",X"00",X"99",X"EE",X"05",X"00",
		X"FF",X"95",X"A0",X"00",X"99",X"F9",X"AA",X"00",X"D9",X"9F",X"AA",X"00",X"00",X"E9",X"99",X"00",
		X"00",X"EE",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"00",X"00",
		X"59",X"00",X"00",X"00",X"59",X"A0",X"00",X"00",X"59",X"EE",X"00",X"00",X"53",X"AA",X"00",X"00",
		X"39",X"EE",X"99",X"00",X"99",X"AA",X"AE",X"EE",X"9F",X"99",X"9A",X"E5",X"FF",X"A9",X"AF",X"99",
		X"99",X"79",X"9A",X"9A",X"99",X"A9",X"99",X"FF",X"FF",X"A9",X"A7",X"A9",X"99",X"9F",X"EA",X"99",
		X"99",X"9F",X"AE",X"A7",X"FF",X"FF",X"EA",X"EA",X"99",X"F9",X"AE",X"AE",X"99",X"99",X"EE",X"EA",
		X"F9",X"99",X"EE",X"AE",X"FF",X"F9",X"5E",X"EA",X"99",X"F9",X"EE",X"AE",X"99",X"FF",X"5E",X"AE",
		X"9E",X"9F",X"E5",X"EA",X"EE",X"F9",X"65",X"AE",X"E5",X"99",X"A5",X"EA",X"EE",X"99",X"DA",X"5E",
		X"AE",X"BE",X"FD",X"A5",X"00",X"AE",X"DD",X"DA",X"00",X"EE",X"AD",X"DD",X"00",X"E0",X"EA",X"DD",
		X"00",X"00",X"0E",X"AD",X"00",X"00",X"00",X"5A",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",X"0E",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"E9",X"90",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"EE",
		X"EE",X"AE",X"99",X"E5",X"EE",X"9A",X"EA",X"99",X"AE",X"A9",X"A9",X"A9",X"AA",X"9A",X"FA",X"9A",
		X"99",X"99",X"A9",X"A9",X"9F",X"99",X"99",X"99",X"FF",X"F9",X"A7",X"A7",X"99",X"F9",X"EA",X"EA",
		X"9F",X"F9",X"AE",X"AE",X"9F",X"9A",X"EA",X"EA",X"FF",X"9A",X"AE",X"AE",X"9F",X"9A",X"EE",X"EA",
		X"9F",X"9A",X"EE",X"AE",X"FF",X"9A",X"EE",X"EA",X"9F",X"9A",X"E5",X"AE",X"9F",X"99",X"EE",X"EA",
		X"99",X"F9",X"5E",X"AE",X"FF",X"F9",X"55",X"55",X"9F",X"F9",X"AA",X"AA",X"99",X"99",X"DD",X"DD",
		X"9E",X"99",X"FD",X"DD",X"EE",X"BE",X"DD",X"DD",X"E5",X"AE",X"AA",X"AA",X"EE",X"EE",X"EE",X"5E",
		X"AE",X"E9",X"90",X"EE",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"A9",X"00",X"00",X"00",X"09",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9F",X"99",X"00",X"00",X"9F",X"EE",X"99",X"00",
		X"9E",X"AA",X"EA",X"00",X"44",X"A9",X"EE",X"9E",X"96",X"99",X"95",X"AA",X"99",X"99",X"95",X"99",
		X"9A",X"04",X"39",X"99",X"99",X"49",X"39",X"99",X"9A",X"A9",X"E9",X"99",X"9A",X"99",X"99",X"A3",
		X"9A",X"49",X"99",X"EA",X"9A",X"9A",X"99",X"EE",X"9A",X"4A",X"99",X"EA",X"E4",X"A9",X"99",X"EA",
		X"9E",X"AA",X"99",X"AE",X"09",X"99",X"99",X"EA",X"99",X"44",X"99",X"AE",X"E9",X"EE",X"99",X"E9",
		X"F9",X"99",X"99",X"33",X"99",X"99",X"99",X"BA",X"99",X"AA",X"F5",X"93",X"99",X"AA",X"55",X"99",
		X"00",X"99",X"EE",X"55",X"00",X"00",X"EA",X"9E",X"00",X"00",X"99",X"99",X"00",X"00",X"00",X"E9",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E3",X"00",X"00",X"00",
		X"9E",X"00",X"00",X"00",X"93",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"EE",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"39",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"E9",X"00",X"00",X"99",X"99",X"00",X"00",X"EA",X"9E",X"00",X"99",X"EE",X"55",
		X"99",X"EE",X"55",X"99",X"99",X"AA",X"F5",X"93",X"99",X"99",X"99",X"BA",X"F9",X"99",X"99",X"33",
		X"E9",X"EE",X"99",X"E9",X"99",X"44",X"99",X"AE",X"09",X"99",X"99",X"EA",X"9E",X"AA",X"99",X"AE",
		X"E4",X"A9",X"99",X"EA",X"9A",X"4A",X"99",X"EA",X"9A",X"9A",X"99",X"EE",X"9A",X"49",X"99",X"EA",
		X"9A",X"99",X"99",X"A3",X"9A",X"A9",X"E9",X"99",X"99",X"49",X"39",X"99",X"9A",X"04",X"39",X"99",
		X"99",X"99",X"95",X"99",X"96",X"99",X"95",X"AA",X"44",X"A9",X"EE",X"9E",X"9E",X"AA",X"EA",X"00",
		X"9F",X"AE",X"99",X"00",X"9F",X"99",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",
		X"E9",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"9A",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"EE",X"00",X"00",X"00",
		X"AA",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"93",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"99",X"00",X"90",X"09",X"99",X"09",X"09",X"22",X"22",X"99",X"99",X"92",X"22",
		X"99",X"99",X"92",X"22",X"21",X"33",X"92",X"22",X"13",X"A3",X"92",X"22",X"71",X"AA",X"92",X"22",
		X"13",X"FF",X"92",X"22",X"22",X"22",X"92",X"22",X"29",X"27",X"92",X"22",X"37",X"44",X"92",X"22",
		X"71",X"46",X"92",X"22",X"11",X"74",X"92",X"22",X"11",X"66",X"92",X"22",X"11",X"66",X"92",X"22",
		X"99",X"66",X"92",X"22",X"77",X"66",X"92",X"22",X"14",X"74",X"92",X"22",X"11",X"76",X"92",X"22",
		X"74",X"74",X"92",X"22",X"37",X"77",X"92",X"22",X"39",X"27",X"92",X"22",X"D3",X"22",X"92",X"22",
		X"13",X"FF",X"92",X"22",X"71",X"22",X"92",X"22",X"13",X"A2",X"92",X"22",X"21",X"33",X"92",X"22",
		X"99",X"00",X"92",X"22",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"05",X"51",X"00",X"00",X"55",X"51",X"50",
		X"00",X"55",X"11",X"55",X"00",X"55",X"11",X"55",X"05",X"55",X"11",X"33",X"55",X"53",X"11",X"33",
		X"55",X"34",X"11",X"73",X"91",X"43",X"99",X"34",X"94",X"93",X"BB",X"35",X"55",X"33",X"BB",X"99",
		X"F1",X"33",X"B9",X"9F",X"11",X"35",X"99",X"99",X"11",X"55",X"95",X"99",X"11",X"55",X"95",X"99",
		X"11",X"55",X"95",X"99",X"11",X"55",X"95",X"99",X"11",X"35",X"B9",X"99",X"31",X"33",X"B9",X"95",
		X"55",X"FF",X"BB",X"99",X"94",X"FF",X"BB",X"31",X"91",X"11",X"FF",X"54",X"55",X"54",X"11",X"1F",
		X"F5",X"55",X"11",X"55",X"0F",X"55",X"11",X"55",X"00",X"55",X"11",X"FF",X"00",X"FF",X"11",X"F0",
		X"00",X"FF",X"51",X"00",X"00",X"0F",X"F1",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"99",X"00",X"00",X"99",X"99",X"00",X"00",X"9F",X"FF",X"00",X"00",
		X"F3",X"33",X"00",X"00",X"F5",X"55",X"00",X"00",X"11",X"59",X"00",X"00",X"11",X"11",X"00",X"00",
		X"99",X"99",X"00",X"00",X"FF",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",
		X"F9",X"FF",X"00",X"00",X"F9",X"FF",X"00",X"00",X"FF",X"FF",X"00",X"00",X"99",X"99",X"00",X"00",
		X"14",X"11",X"00",X"00",X"11",X"FF",X"00",X"00",X"9F",X"F5",X"00",X"00",X"9E",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"F9",X"99",X"00",X"00",X"0F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"99",X"99",X"00",X"00",X"EE",X"90",X"00",X"00",X"EE",X"09",X"00",X"00",X"29",X"90",X"00",X"00",
		X"22",X"09",X"00",X"00",X"22",X"90",X"00",X"00",X"22",X"90",X"00",X"00",X"99",X"09",X"00",X"00",
		X"99",X"99",X"00",X"00",X"22",X"F3",X"09",X"00",X"22",X"33",X"90",X"00",X"22",X"99",X"90",X"00",
		X"99",X"99",X"99",X"00",X"33",X"3F",X"99",X"00",X"23",X"33",X"9F",X"00",X"99",X"99",X"FF",X"00",
		X"22",X"92",X"F9",X"00",X"22",X"92",X"F9",X"00",X"22",X"92",X"39",X"00",X"22",X"92",X"99",X"00",
		X"29",X"99",X"9F",X"00",X"22",X"22",X"FF",X"00",X"22",X"22",X"F9",X"00",X"22",X"22",X"F0",X"00",
		X"22",X"29",X"F9",X"00",X"22",X"29",X"90",X"00",X"92",X"29",X"00",X"00",X"22",X"22",X"00",X"00",
		X"22",X"29",X"09",X"00",X"22",X"29",X"90",X"00",X"22",X"29",X"00",X"00",X"22",X"29",X"09",X"00",
		X"11",X"19",X"09",X"00",X"11",X"19",X"00",X"00",X"11",X"19",X"90",X"00",X"11",X"19",X"09",X"00",
		X"11",X"12",X"00",X"00",X"11",X"12",X"00",X"00",X"11",X"19",X"90",X"00",X"22",X"29",X"F9",X"00",
		X"22",X"11",X"F0",X"00",X"99",X"11",X"F9",X"00",X"11",X"11",X"FF",X"00",X"11",X"99",X"9F",X"00",
		X"11",X"92",X"99",X"00",X"11",X"92",X"39",X"00",X"11",X"92",X"F9",X"00",X"22",X"92",X"F9",X"00",
		X"99",X"99",X"FF",X"00",X"13",X"33",X"9F",X"00",X"33",X"3F",X"99",X"00",X"99",X"99",X"99",X"00",
		X"22",X"99",X"90",X"00",X"22",X"33",X"90",X"00",X"22",X"F3",X"09",X"00",X"99",X"99",X"00",X"00",
		X"99",X"09",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"90",X"00",X"00",X"11",X"09",X"00",X"00",
		X"19",X"90",X"00",X"00",X"EE",X"09",X"00",X"00",X"EE",X"90",X"00",X"00",X"99",X"99",X"00",X"00",
		X"91",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"59",X"50",X"00",X"00",X"55",X"55",X"00",X"00",
		X"5F",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"11",X"55",X"00",X"00",X"1F",X"55",X"00",X"00",
		X"15",X"15",X"50",X"00",X"11",X"11",X"55",X"00",X"11",X"11",X"55",X"00",X"F1",X"51",X"55",X"00",
		X"11",X"33",X"55",X"00",X"11",X"33",X"55",X"00",X"11",X"53",X"55",X"00",X"11",X"55",X"11",X"00",
		X"11",X"55",X"11",X"00",X"51",X"F9",X"11",X"10",X"51",X"99",X"11",X"99",X"55",X"99",X"11",X"90",
		X"55",X"9B",X"19",X"09",X"55",X"B9",X"11",X"09",X"55",X"B9",X"F1",X"99",X"55",X"B9",X"BF",X"90",
		X"55",X"BB",X"BB",X"99",X"F5",X"9B",X"9B",X"09",X"F5",X"FB",X"99",X"09",X"05",X"1F",X"9D",X"09",
		X"0F",X"91",X"DD",X"00",X"00",X"91",X"D9",X"00",X"00",X"99",X"99",X"59",X"00",X"95",X"99",X"55",
		X"99",X"99",X"12",X"99",X"99",X"99",X"91",X"99",X"99",X"19",X"99",X"99",X"99",X"12",X"93",X"F9",
		X"99",X"55",X"FF",X"00",X"90",X"55",X"99",X"99",X"90",X"00",X"9F",X"99",X"00",X"99",X"F9",X"FF",
		X"90",X"99",X"99",X"00",X"09",X"00",X"9F",X"F0",X"00",X"09",X"F9",X"F0",X"00",X"09",X"39",X"1F",
		X"00",X"00",X"19",X"11",X"00",X"00",X"12",X"99",X"00",X"00",X"F1",X"90",X"00",X"00",X"F1",X"99",
		X"00",X"00",X"9F",X"09",X"00",X"00",X"9F",X"00",X"00",X"00",X"90",X"90",X"00",X"00",X"90",X"00",
		X"00",X"00",X"90",X"00",X"00",X"00",X"99",X"90",X"00",X"00",X"99",X"90",X"00",X"00",X"06",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"09",X"00",X"09",X"00",X"13",X"99",X"90",X"00",X"91",X"33",X"09",X"00",X"99",X"5F",X"99",X"90",
		X"19",X"55",X"33",X"00",X"11",X"55",X"FF",X"09",X"55",X"15",X"5F",X"90",X"F5",X"11",X"5F",X"99",
		X"FF",X"11",X"55",X"99",X"FF",X"F1",X"55",X"11",X"FF",X"5F",X"55",X"11",X"1F",X"59",X"11",X"19",
		X"11",X"99",X"11",X"99",X"11",X"99",X"11",X"99",X"51",X"95",X"BF",X"93",X"55",X"95",X"BB",X"55",
		X"55",X"F9",X"99",X"F5",X"55",X"F9",X"99",X"55",X"F5",X"FF",X"99",X"15",X"FF",X"1F",X"99",X"11",
		X"0F",X"11",X"99",X"91",X"0F",X"11",X"99",X"F1",X"00",X"51",X"B9",X"FF",X"00",X"F5",X"FB",X"F9",
		X"00",X"55",X"11",X"F9",X"00",X"F5",X"11",X"99",X"00",X"F5",X"99",X"99",X"00",X"F5",X"99",X"19",
		X"00",X"FF",X"99",X"11",X"00",X"FF",X"99",X"91",X"00",X"FF",X"99",X"95",X"00",X"0F",X"99",X"95",
		X"55",X"F3",X"00",X"00",X"55",X"FF",X"90",X"00",X"11",X"F1",X"90",X"00",X"11",X"11",X"00",X"00",
		X"11",X"11",X"00",X"00",X"9F",X"11",X"90",X"00",X"F5",X"11",X"09",X"00",X"99",X"19",X"00",X"00",
		X"9B",X"19",X"09",X"00",X"9B",X"19",X"99",X"00",X"BB",X"B1",X"99",X"00",X"BB",X"9B",X"39",X"00",
		X"B9",X"99",X"99",X"00",X"BB",X"29",X"FF",X"00",X"BB",X"29",X"F3",X"00",X"1F",X"9D",X"F3",X"99",
		X"11",X"9D",X"FF",X"FF",X"11",X"DD",X"99",X"90",X"11",X"DF",X"91",X"F9",X"11",X"D9",X"F9",X"0F",
		X"11",X"11",X"98",X"90",X"11",X"55",X"98",X"F9",X"11",X"55",X"8F",X"FF",X"21",X"FF",X"89",X"1F",
		X"F1",X"FF",X"11",X"5F",X"F1",X"00",X"F1",X"F3",X"F1",X"00",X"0F",X"33",X"01",X"00",X"00",X"33",
		X"00",X"00",X"90",X"33",X"00",X"00",X"99",X"39",X"00",X"00",X"F9",X"39",X"00",X"00",X"FF",X"00",
		X"00",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"9C",X"99",X"99",X"00",X"C9",X"99",X"99",X"00",
		X"65",X"99",X"99",X"00",X"65",X"EB",X"99",X"90",X"65",X"CA",X"C9",X"99",X"99",X"AA",X"0C",X"99",
		X"A9",X"EA",X"EC",X"C9",X"EE",X"BB",X"AB",X"B9",X"EB",X"BE",X"BA",X"BC",X"EB",X"BB",X"EE",X"9B",
		X"5E",X"BB",X"BB",X"CB",X"E5",X"EB",X"BB",X"9C",X"EB",X"FE",X"BB",X"BC",X"EB",X"B5",X"5B",X"BC",
		X"6F",X"BA",X"BB",X"9C",X"B6",X"BA",X"BB",X"BC",X"9B",X"BA",X"B5",X"EC",X"9C",X"BA",X"BB",X"BC",
		X"5C",X"BA",X"5B",X"EC",X"BC",X"BB",X"BB",X"BC",X"B6",X"FB",X"FB",X"9C",X"BB",X"CB",X"BB",X"C9",
		X"CC",X"CC",X"FB",X"5F",X"00",X"99",X"BB",X"09",X"00",X"00",X"CC",X"C9",X"00",X"00",X"99",X"C9",
		X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",
		X"00",X"90",X"99",X"90",X"00",X"99",X"99",X"C9",X"09",X"99",X"CC",X"C9",X"00",X"99",X"AB",X"09",
		X"90",X"CC",X"BA",X"5F",X"00",X"CA",X"AB",X"C9",X"B6",X"AA",X"BB",X"9C",X"BC",X"AA",X"BB",X"BC",
		X"5C",X"BA",X"BB",X"EC",X"9C",X"AA",X"BB",X"BC",X"9B",X"BA",X"BB",X"EC",X"BA",X"BA",X"BB",X"BC",
		X"AA",X"BA",X"BB",X"9C",X"EB",X"BE",X"5B",X"BC",X"EB",X"EF",X"BB",X"BC",X"EE",X"FB",X"BB",X"9C",
		X"55",X"BB",X"BB",X"CB",X"EB",X"BB",X"55",X"9B",X"EB",X"BE",X"BF",X"BC",X"EE",X"BB",X"FB",X"B9",
		X"A9",X"FB",X"EC",X"CA",X"99",X"6B",X"0A",X"A0",X"65",X"BB",X"C9",X"00",X"65",X"EB",X"A0",X"00",
		X"65",X"9A",X"00",X"00",X"C9",X"A0",X"00",X"00",X"9C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"D9",X"00",X"00",X"D9",X"99",X"00",X"00",X"99",X"99",
		X"00",X"D9",X"99",X"FF",X"0D",X"5A",X"99",X"99",X"09",X"EA",X"99",X"99",X"D9",X"AE",X"9E",X"99",
		X"59",X"EE",X"9E",X"99",X"99",X"AE",X"E5",X"99",X"93",X"E9",X"EE",X"99",X"93",X"99",X"AA",X"9E",
		X"9A",X"EE",X"AA",X"99",X"A3",X"EE",X"AA",X"99",X"99",X"EF",X"AA",X"99",X"9F",X"FF",X"A5",X"99",
		X"59",X"FF",X"55",X"59",X"59",X"FF",X"99",X"59",X"59",X"FF",X"99",X"59",X"59",X"AF",X"AA",X"59",
		X"59",X"AA",X"AA",X"F9",X"59",X"3A",X"7A",X"33",X"59",X"93",X"53",X"A3",X"09",X"99",X"3A",X"99",
		X"F3",X"55",X"99",X"99",X"FF",X"EE",X"99",X"99",X"F0",X"EE",X"99",X"AA",X"F0",X"EA",X"99",X"00",
		X"FF",X"E7",X"AA",X"00",X"FF",X"E9",X"00",X"00",X"0F",X"AA",X"00",X"00",X"0F",X"A0",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"99",X"99",X"00",X"00",X"E0",X"99",X"00",X"00",X"EE",X"99",X"00",
		X"00",X"E9",X"99",X"00",X"D9",X"9F",X"AA",X"00",X"99",X"F9",X"AA",X"00",X"FF",X"95",X"A0",X"00",
		X"99",X"EE",X"05",X"00",X"EE",X"AA",X"99",X"00",X"EE",X"AA",X"99",X"00",X"AE",X"AA",X"99",X"00",
		X"AE",X"AA",X"F9",X"00",X"AA",X"AA",X"F9",X"00",X"AA",X"9A",X"F9",X"00",X"AA",X"AA",X"F9",X"00",
		X"AA",X"9A",X"F9",X"00",X"AA",X"AA",X"F9",X"00",X"AA",X"AA",X"F9",X"00",X"AA",X"AA",X"99",X"00",
		X"AA",X"94",X"99",X"F0",X"AA",X"AA",X"99",X"F0",X"AA",X"AA",X"9A",X"F0",X"AA",X"A7",X"99",X"F0",
		X"AA",X"99",X"99",X"00",X"A9",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"99",X"3A",X"00",X"00",
		X"99",X"99",X"90",X"00",X"99",X"09",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"09",X"09",X"00",X"00",X"92",X"99",X"00",X"00",X"2D",X"99",X"09",X"90",
		X"F2",X"22",X"92",X"99",X"67",X"22",X"22",X"99",X"27",X"11",X"22",X"22",X"21",X"11",X"99",X"22",
		X"11",X"99",X"39",X"22",X"1E",X"99",X"13",X"99",X"19",X"99",X"71",X"91",X"19",X"99",X"77",X"11",
		X"19",X"99",X"77",X"09",X"19",X"99",X"77",X"13",X"19",X"99",X"77",X"13",X"17",X"99",X"77",X"13",
		X"DF",X"93",X"77",X"33",X"ED",X"9F",X"77",X"33",X"1E",X"F3",X"77",X"33",X"11",X"99",X"77",X"33",
		X"71",X"99",X"75",X"33",X"57",X"99",X"F7",X"33",X"2F",X"77",X"11",X"99",X"02",X"2A",X"33",X"11",
		X"09",X"22",X"99",X"19",X"00",X"00",X"22",X"91",X"00",X"00",X"52",X"21",X"00",X"00",X"22",X"21",
		X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"92",X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"22",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"1A",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"09",X"00",X"00",X"00",X"09",X"00",X"00",X"99",X"92",X"00",X"00",X"99",X"22",
		X"00",X"00",X"22",X"21",X"00",X"09",X"22",X"21",X"00",X"99",X"22",X"91",X"09",X"22",X"99",X"19",
		X"92",X"2A",X"33",X"11",X"24",X"77",X"11",X"99",X"47",X"99",X"77",X"33",X"71",X"99",X"DD",X"33",
		X"11",X"99",X"77",X"33",X"1E",X"99",X"77",X"33",X"ED",X"99",X"77",X"33",X"DF",X"93",X"77",X"33",
		X"17",X"99",X"77",X"13",X"19",X"99",X"77",X"13",X"19",X"99",X"77",X"13",X"19",X"99",X"77",X"09",
		X"19",X"99",X"75",X"11",X"19",X"9F",X"71",X"91",X"1E",X"F9",X"13",X"99",X"11",X"99",X"39",X"22",
		X"21",X"11",X"99",X"22",X"27",X"11",X"22",X"22",X"67",X"22",X"55",X"00",X"F2",X"22",X"02",X"00",
		X"2D",X"99",X"00",X"00",X"92",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",X"29",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"72",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",X"12",X"00",X"00",X"00",
		X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"15",X"00",X"00",X"00",
		X"15",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"22",X"00",X"00",X"00",
		X"29",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0F",X"00",X"00",X"00",X"0F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"9F",X"00",X"00",X"00",X"5F",X"00",X"00",X"00",X"9F",X"00",X"00",
		X"00",X"5F",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"AF",X"00",X"00",X"00",X"AA",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"55",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"9A",X"9A",X"9A",X"00",X"AB",X"AB",X"AB",X"00",X"BD",X"BD",X"BD",X"00",X"BB",X"BB",X"BB",
		X"00",X"5B",X"5B",X"5B",X"00",X"BA",X"BA",X"BA",X"00",X"DD",X"99",X"99",X"00",X"99",X"99",X"99",
		X"09",X"DE",X"EE",X"55",X"9D",X"99",X"B5",X"99",X"DD",X"DE",X"5B",X"EE",X"99",X"EE",X"B5",X"99",
		X"DD",X"E9",X"99",X"AB",X"99",X"E9",X"FE",X"BA",X"DD",X"99",X"F9",X"AB",X"99",X"EE",X"F5",X"BA",
		X"AA",X"BB",X"F5",X"AB",X"AB",X"99",X"F9",X"BA",X"BA",X"59",X"F5",X"AB",X"AB",X"B9",X"B5",X"9A",
		X"BA",X"5B",X"5B",X"99",X"AB",X"A5",X"55",X"FF",X"BA",X"BB",X"5B",X"99",X"0B",X"A5",X"F5",X"55",
		X"00",X"BA",X"99",X"95",X"00",X"AB",X"99",X"99",X"00",X"99",X"99",X"99",X"00",X"BA",X"BA",X"BA",
		X"00",X"AB",X"AB",X"AB",X"00",X"BB",X"BB",X"BB",X"00",X"B5",X"B5",X"B5",X"00",X"AB",X"AB",X"AB",
		X"99",X"99",X"90",X"00",X"AB",X"A9",X"A0",X"00",X"BD",X"BD",X"99",X"00",X"BB",X"B9",X"9D",X"00",
		X"59",X"5B",X"59",X"00",X"BA",X"B9",X"B9",X"00",X"9D",X"DD",X"99",X"00",X"99",X"DD",X"99",X"00",
		X"EE",X"BB",X"99",X"00",X"9E",X"DD",X"99",X"00",X"E9",X"BB",X"99",X"00",X"AE",X"DD",X"99",X"00",
		X"E9",X"BB",X"99",X"00",X"A9",X"BB",X"99",X"00",X"99",X"BB",X"99",X"00",X"A9",X"BB",X"99",X"00",
		X"99",X"AB",X"99",X"00",X"A9",X"BB",X"99",X"00",X"99",X"AB",X"99",X"00",X"A9",X"BB",X"99",X"00",
		X"99",X"AA",X"99",X"00",X"99",X"BB",X"99",X"00",X"99",X"AA",X"99",X"00",X"99",X"B9",X"99",X"00",
		X"59",X"AA",X"99",X"00",X"55",X"B9",X"99",X"00",X"99",X"99",X"99",X"00",X"AB",X"A9",X"9A",X"00",
		X"BA",X"BA",X"9A",X"00",X"BB",X"B9",X"9A",X"00",X"B5",X"B5",X"90",X"00",X"AB",X"A9",X"90",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"B0",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BF",X"BB",X"00",X"00",X"BF",X"BB",X"00",X"00",X"BF",X"BB",X"BB",X"00",X"BF",X"BB",X"BB",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BF",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"BF",X"BB",
		X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"BF",X"00",X"BB",X"0B",
		X"BF",X"00",X"BB",X"00",X"BF",X"00",X"BF",X"B0",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",
		X"BF",X"00",X"0B",X"BB",X"BF",X"00",X"0B",X"BB",X"BF",X"00",X"0B",X"BB",X"BF",X"00",X"0B",X"BB",
		X"BF",X"00",X"0B",X"BB",X"BF",X"00",X"0B",X"BB",X"BF",X"00",X"0B",X"BB",X"BF",X"BB",X"0B",X"BB",
		X"BF",X"BB",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",X"0B",X"BB",X"0B",X"BB",X"00",X"FB",X"0B",X"BB",
		X"00",X"BB",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"FB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"B0",
		X"0B",X"BB",X"BB",X"B0",X"BB",X"FB",X"BB",X"B0",X"BB",X"BB",X"BF",X"B0",X"BB",X"B0",X"BB",X"B0",
		X"BB",X"00",X"00",X"B0",X"BF",X"00",X"00",X"B0",X"BB",X"00",X"00",X"B0",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",
		X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"FF",X"00",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"FB",X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",
		X"BB",X"00",X"BB",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"FB",X"0B",
		X"BB",X"00",X"BB",X"00",X"BB",X"00",X"BB",X"B0",X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",
		X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",
		X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",
		X"BB",X"FB",X"0B",X"BB",X"BB",X"BF",X"0B",X"BB",X"0B",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",
		X"00",X"BB",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"BF",X"BB",
		X"0B",X"BB",X"BB",X"FB",X"BB",X"BB",X"BB",X"FB",X"FB",X"BB",X"BB",X"FB",X"BB",X"B0",X"BB",X"FB",
		X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",X"00",X"00",
		X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"FF",X"BB",X"00",X"BB",X"BB",X"BB",X"00",
		X"BB",X"BB",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",X"BB",X"BB",X"00",X"BB",X"BB",
		X"BB",X"00",X"BB",X"BB",X"BF",X"00",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"BF",X"00",X"BB",X"0B",
		X"BF",X"00",X"FB",X"00",X"BF",X"00",X"BF",X"B0",X"BF",X"00",X"BB",X"BB",X"BF",X"00",X"FB",X"BB",
		X"BF",X"00",X"0F",X"BB",X"BF",X"00",X"0F",X"BB",X"BF",X"00",X"0B",X"BB",X"BF",X"00",X"0B",X"BB",
		X"BF",X"00",X"0B",X"BB",X"BF",X"00",X"0B",X"BB",X"BB",X"00",X"0B",X"BB",X"BB",X"BB",X"0B",X"BB",
		X"BB",X"FB",X"0B",X"BB",X"BB",X"BF",X"0B",X"BB",X"0B",X"BB",X"0B",X"BB",X"00",X"BB",X"0B",X"BB",
		X"00",X"BB",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",
		X"FF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",
		X"00",X"FF",X"00",X"00",X"00",X"FF",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"BB",X"BB",X"BB",
		X"0B",X"BB",X"FF",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BB",X"BF",X"B0",X"BB",X"BB",
		X"BF",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"B0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BF",X"BB",X"00",X"00",
		X"FF",X"BF",X"00",X"00",X"FF",X"BB",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",
		X"FF",X"BB",X"00",X"00",X"FF",X"BB",X"00",X"00",X"FF",X"BB",X"BB",X"00",X"FF",X"BB",X"BB",X"00",
		X"BB",X"FF",X"BB",X"BB",X"BB",X"FF",X"BB",X"BB",X"00",X"BB",X"FF",X"BB",X"BB",X"00",X"BF",X"BB",
		X"BB",X"00",X"BB",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"BB",X"BB",X"FF",X"00",X"BB",X"0B",
		X"FF",X"00",X"BB",X"00",X"FF",X"00",X"BF",X"B0",X"FB",X"00",X"FF",X"BB",X"FB",X"00",X"BB",X"BB",
		X"FF",X"00",X"0B",X"BB",X"FF",X"00",X"0B",X"BB",X"FF",X"00",X"0B",X"BB",X"FF",X"00",X"0B",X"BB",
		X"FF",X"00",X"0B",X"BB",X"FF",X"00",X"0B",X"BB",X"FF",X"00",X"0B",X"BB",X"FF",X"BB",X"0B",X"BB",
		X"FF",X"BB",X"0B",X"BB",X"BF",X"BB",X"0B",X"BB",X"0B",X"FB",X"0B",X"BB",X"00",X"FF",X"0B",X"BB",
		X"00",X"BB",X"0B",X"BB",X"00",X"00",X"0B",X"BB",X"00",X"00",X"00",X"FB",X"00",X"00",X"00",X"BB",
		X"BF",X"00",X"00",X"00",X"BF",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"0B",X"B0",X"00",X"00",
		X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",X"00",X"BB",X"00",X"00",
		X"00",X"FB",X"00",X"00",X"00",X"BF",X"BB",X"00",X"00",X"BB",X"BB",X"00",X"00",X"BB",X"BB",X"BB",
		X"0B",X"BF",X"BB",X"BB",X"BB",X"FF",X"FF",X"BB",X"BB",X"FB",X"FF",X"BB",X"BB",X"B0",X"BB",X"BB",
		X"BB",X"00",X"00",X"BB",X"BF",X"00",X"00",X"BB",X"FF",X"00",X"00",X"BB",X"F0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"0B",X"00",X"00",X"00",X"BB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",
		X"FB",X"BB",X"00",X"00",X"FB",X"BB",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"11",
		X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"11",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"00",X"00",
		X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"11",X"00",X"00",X"01",X"11",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"11",
		X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"00",X"00",X"00",X"11",
		X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",X"10",X"11",X"11",X"11",X"10",X"11",X"11",X"11",
		X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"10",X"11",X"11",X"11",X"10",X"11",X"11",X"11",
		X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"10",X"11",X"11",X"11",X"10",X"11",X"11",X"11",
		X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"10",X"00",X"00",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"11",X"10",X"11",X"11",X"11",X"10",X"11",
		X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",X"10",X"11",X"11",X"11",X"10",X"11",X"11",X"10",
		X"10",X"00",X"11",X"00",X"10",X"00",X"10",X"00",X"10",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"10",X"00",X"01",X"00",X"10",X"00",X"11",X"00",X"10",X"11",X"11",X"11",X"10",X"11",X"11",X"11",
		X"10",X"00",X"00",X"11",X"10",X"00",X"00",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"11",
		X"11",X"00",X"10",X"11",X"11",X"00",X"10",X"11",X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",
		X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",X"10",X"00",X"10",X"11",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"0A",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",
		X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"0E",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"A0",X"00",
		X"00",X"00",X"A0",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"AA",X"00",X"00",X"00",X"00",X"00",
		X"00",X"0E",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"55",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"0B",X"99",X"00",
		X"00",X"FF",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"09",X"00",X"99",X"09",X"99",X"00",X"99",X"99",X"99",
		X"99",X"99",X"99",X"F5",X"EE",X"EE",X"EE",X"EE",X"BB",X"BB",X"BB",X"BB",X"44",X"45",X"99",X"5F",
		X"77",X"77",X"99",X"99",X"33",X"59",X"55",X"9B",X"55",X"53",X"FF",X"B5",X"5F",X"39",X"FF",X"99",
		X"FE",X"99",X"FF",X"99",X"99",X"99",X"FF",X"99",X"59",X"93",X"FF",X"99",X"59",X"93",X"FF",X"99",
		X"59",X"93",X"FF",X"99",X"59",X"93",X"FF",X"99",X"99",X"93",X"FF",X"99",X"FF",X"93",X"FF",X"99",
		X"55",X"93",X"FF",X"99",X"55",X"59",X"FF",X"55",X"33",X"59",X"55",X"95",X"77",X"77",X"99",X"99",
		X"F4",X"45",X"99",X"55",X"BF",X"BB",X"BB",X"BB",X"EF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"F5",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"90",X"00",X"00",X"00",X"90",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"E9",X"00",X"00",X"00",X"BE",X"00",X"00",X"00",
		X"E1",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"91",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",
		X"9E",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",X"99",X"00",X"00",X"00",
		X"9E",X"00",X"00",X"00",X"9E",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",X"E1",X"00",X"00",X"00",
		X"BF",X"00",X"00",X"00",X"E0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
